`timescale 1ns / 1ps
`include "param.v"

module systolic_loader_p (
CLK,
    i_Psram_Addr,
    i_Psram_En,
    i_Psram_Valid_1buf,
    o_Psram_Addr_To_Sram,
    o_Psram_En_To_Sram,
    o_Psram_Valid_To_Systolic );

    input CLK;
    input [`BIT_ADDR-1:0] i_Psram_Addr;
    input [`PE_COL-1:0] i_Psram_En;
    input [`PE_COL-1:0] i_Psram_Valid_1buf;
    output [`BIT_ADDR*`PE_COL-1:0] o_Psram_Addr_To_Sram;
    output [`PE_COL-1:0] o_Psram_En_To_Sram;
    output [`PE_COL-1:0] o_Psram_Valid_To_Systolic;

    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_1 [0:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_2 [1:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_3 [2:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_4 [3:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_5 [4:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_6 [5:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_7 [6:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_8 [7:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_9 [8:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_10 [9:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_11 [10:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_12 [11:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_13 [12:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_14 [13:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_15 [14:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_16 [15:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_17 [16:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_18 [17:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_19 [18:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_20 [19:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_21 [20:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_22 [21:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_23 [22:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_24 [23:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_25 [24:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_26 [25:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_27 [26:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_28 [27:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_29 [28:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_30 [29:0];
    reg [`BIT_ADDR-1:0] Psram_Addr_To_Sram_FIFO_31 [30:0];
    reg  Psram_En_To_Sram_FIFO_1 [0:0];
    reg  Psram_En_To_Sram_FIFO_2 [1:0];
    reg  Psram_En_To_Sram_FIFO_3 [2:0];
    reg  Psram_En_To_Sram_FIFO_4 [3:0];
    reg  Psram_En_To_Sram_FIFO_5 [4:0];
    reg  Psram_En_To_Sram_FIFO_6 [5:0];
    reg  Psram_En_To_Sram_FIFO_7 [6:0];
    reg  Psram_En_To_Sram_FIFO_8 [7:0];
    reg  Psram_En_To_Sram_FIFO_9 [8:0];
    reg  Psram_En_To_Sram_FIFO_10 [9:0];
    reg  Psram_En_To_Sram_FIFO_11 [10:0];
    reg  Psram_En_To_Sram_FIFO_12 [11:0];
    reg  Psram_En_To_Sram_FIFO_13 [12:0];
    reg  Psram_En_To_Sram_FIFO_14 [13:0];
    reg  Psram_En_To_Sram_FIFO_15 [14:0];
    reg  Psram_En_To_Sram_FIFO_16 [15:0];
    reg  Psram_En_To_Sram_FIFO_17 [16:0];
    reg  Psram_En_To_Sram_FIFO_18 [17:0];
    reg  Psram_En_To_Sram_FIFO_19 [18:0];
    reg  Psram_En_To_Sram_FIFO_20 [19:0];
    reg  Psram_En_To_Sram_FIFO_21 [20:0];
    reg  Psram_En_To_Sram_FIFO_22 [21:0];
    reg  Psram_En_To_Sram_FIFO_23 [22:0];
    reg  Psram_En_To_Sram_FIFO_24 [23:0];
    reg  Psram_En_To_Sram_FIFO_25 [24:0];
    reg  Psram_En_To_Sram_FIFO_26 [25:0];
    reg  Psram_En_To_Sram_FIFO_27 [26:0];
    reg  Psram_En_To_Sram_FIFO_28 [27:0];
    reg  Psram_En_To_Sram_FIFO_29 [28:0];
    reg  Psram_En_To_Sram_FIFO_30 [29:0];
    reg  Psram_En_To_Sram_FIFO_31 [30:0];
    reg  Psram_Valid_To_Systolic_FIFO_1 [0:0];
    reg  Psram_Valid_To_Systolic_FIFO_2 [1:0];
    reg  Psram_Valid_To_Systolic_FIFO_3 [2:0];
    reg  Psram_Valid_To_Systolic_FIFO_4 [3:0];
    reg  Psram_Valid_To_Systolic_FIFO_5 [4:0];
    reg  Psram_Valid_To_Systolic_FIFO_6 [5:0];
    reg  Psram_Valid_To_Systolic_FIFO_7 [6:0];
    reg  Psram_Valid_To_Systolic_FIFO_8 [7:0];
    reg  Psram_Valid_To_Systolic_FIFO_9 [8:0];
    reg  Psram_Valid_To_Systolic_FIFO_10 [9:0];
    reg  Psram_Valid_To_Systolic_FIFO_11 [10:0];
    reg  Psram_Valid_To_Systolic_FIFO_12 [11:0];
    reg  Psram_Valid_To_Systolic_FIFO_13 [12:0];
    reg  Psram_Valid_To_Systolic_FIFO_14 [13:0];
    reg  Psram_Valid_To_Systolic_FIFO_15 [14:0];
    reg  Psram_Valid_To_Systolic_FIFO_16 [15:0];
    reg  Psram_Valid_To_Systolic_FIFO_17 [16:0];
    reg  Psram_Valid_To_Systolic_FIFO_18 [17:0];
    reg  Psram_Valid_To_Systolic_FIFO_19 [18:0];
    reg  Psram_Valid_To_Systolic_FIFO_20 [19:0];
    reg  Psram_Valid_To_Systolic_FIFO_21 [20:0];
    reg  Psram_Valid_To_Systolic_FIFO_22 [21:0];
    reg  Psram_Valid_To_Systolic_FIFO_23 [22:0];
    reg  Psram_Valid_To_Systolic_FIFO_24 [23:0];
    reg  Psram_Valid_To_Systolic_FIFO_25 [24:0];
    reg  Psram_Valid_To_Systolic_FIFO_26 [25:0];
    reg  Psram_Valid_To_Systolic_FIFO_27 [26:0];
    reg  Psram_Valid_To_Systolic_FIFO_28 [27:0];
    reg  Psram_Valid_To_Systolic_FIFO_29 [28:0];
    reg  Psram_Valid_To_Systolic_FIFO_30 [29:0];
    reg  Psram_Valid_To_Systolic_FIFO_31 [30:0];
    // Psram_Addr_To_Sram Assignments
    assign o_Psram_Addr_To_Sram[0*`BIT_ADDR +: `BIT_ADDR] = i_Psram_Addr;
    assign o_Psram_Addr_To_Sram[1*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_1[0];
    assign o_Psram_Addr_To_Sram[2*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_2[0];
    assign o_Psram_Addr_To_Sram[3*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_3[0];
    assign o_Psram_Addr_To_Sram[4*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_4[0];
    assign o_Psram_Addr_To_Sram[5*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_5[0];
    assign o_Psram_Addr_To_Sram[6*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_6[0];
    assign o_Psram_Addr_To_Sram[7*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_7[0];
    assign o_Psram_Addr_To_Sram[8*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_8[0];
    assign o_Psram_Addr_To_Sram[9*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_9[0];
    assign o_Psram_Addr_To_Sram[10*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_10[0];
    assign o_Psram_Addr_To_Sram[11*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_11[0];
    assign o_Psram_Addr_To_Sram[12*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_12[0];
    assign o_Psram_Addr_To_Sram[13*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_13[0];
    assign o_Psram_Addr_To_Sram[14*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_14[0];
    assign o_Psram_Addr_To_Sram[15*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_15[0];
    assign o_Psram_Addr_To_Sram[16*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_16[0];
    assign o_Psram_Addr_To_Sram[17*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_17[0];
    assign o_Psram_Addr_To_Sram[18*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_18[0];
    assign o_Psram_Addr_To_Sram[19*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_19[0];
    assign o_Psram_Addr_To_Sram[20*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_20[0];
    assign o_Psram_Addr_To_Sram[21*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_21[0];
    assign o_Psram_Addr_To_Sram[22*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_22[0];
    assign o_Psram_Addr_To_Sram[23*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_23[0];
    assign o_Psram_Addr_To_Sram[24*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_24[0];
    assign o_Psram_Addr_To_Sram[25*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_25[0];
    assign o_Psram_Addr_To_Sram[26*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_26[0];
    assign o_Psram_Addr_To_Sram[27*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_27[0];
    assign o_Psram_Addr_To_Sram[28*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_28[0];
    assign o_Psram_Addr_To_Sram[29*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_29[0];
    assign o_Psram_Addr_To_Sram[30*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_30[0];
    assign o_Psram_Addr_To_Sram[31*`BIT_ADDR +: `BIT_ADDR] = Psram_Addr_To_Sram_FIFO_31[0];

    // Psram_En_To_Sram Assignments
    assign o_Psram_En_To_Sram[0*1 +: 1] = i_Psram_En;
    assign o_Psram_En_To_Sram[1*1 +: 1] = Psram_En_To_Sram_FIFO_1[0];
    assign o_Psram_En_To_Sram[2*1 +: 1] = Psram_En_To_Sram_FIFO_2[0];
    assign o_Psram_En_To_Sram[3*1 +: 1] = Psram_En_To_Sram_FIFO_3[0];
    assign o_Psram_En_To_Sram[4*1 +: 1] = Psram_En_To_Sram_FIFO_4[0];
    assign o_Psram_En_To_Sram[5*1 +: 1] = Psram_En_To_Sram_FIFO_5[0];
    assign o_Psram_En_To_Sram[6*1 +: 1] = Psram_En_To_Sram_FIFO_6[0];
    assign o_Psram_En_To_Sram[7*1 +: 1] = Psram_En_To_Sram_FIFO_7[0];
    assign o_Psram_En_To_Sram[8*1 +: 1] = Psram_En_To_Sram_FIFO_8[0];
    assign o_Psram_En_To_Sram[9*1 +: 1] = Psram_En_To_Sram_FIFO_9[0];
    assign o_Psram_En_To_Sram[10*1 +: 1] = Psram_En_To_Sram_FIFO_10[0];
    assign o_Psram_En_To_Sram[11*1 +: 1] = Psram_En_To_Sram_FIFO_11[0];
    assign o_Psram_En_To_Sram[12*1 +: 1] = Psram_En_To_Sram_FIFO_12[0];
    assign o_Psram_En_To_Sram[13*1 +: 1] = Psram_En_To_Sram_FIFO_13[0];
    assign o_Psram_En_To_Sram[14*1 +: 1] = Psram_En_To_Sram_FIFO_14[0];
    assign o_Psram_En_To_Sram[15*1 +: 1] = Psram_En_To_Sram_FIFO_15[0];
    assign o_Psram_En_To_Sram[16*1 +: 1] = Psram_En_To_Sram_FIFO_16[0];
    assign o_Psram_En_To_Sram[17*1 +: 1] = Psram_En_To_Sram_FIFO_17[0];
    assign o_Psram_En_To_Sram[18*1 +: 1] = Psram_En_To_Sram_FIFO_18[0];
    assign o_Psram_En_To_Sram[19*1 +: 1] = Psram_En_To_Sram_FIFO_19[0];
    assign o_Psram_En_To_Sram[20*1 +: 1] = Psram_En_To_Sram_FIFO_20[0];
    assign o_Psram_En_To_Sram[21*1 +: 1] = Psram_En_To_Sram_FIFO_21[0];
    assign o_Psram_En_To_Sram[22*1 +: 1] = Psram_En_To_Sram_FIFO_22[0];
    assign o_Psram_En_To_Sram[23*1 +: 1] = Psram_En_To_Sram_FIFO_23[0];
    assign o_Psram_En_To_Sram[24*1 +: 1] = Psram_En_To_Sram_FIFO_24[0];
    assign o_Psram_En_To_Sram[25*1 +: 1] = Psram_En_To_Sram_FIFO_25[0];
    assign o_Psram_En_To_Sram[26*1 +: 1] = Psram_En_To_Sram_FIFO_26[0];
    assign o_Psram_En_To_Sram[27*1 +: 1] = Psram_En_To_Sram_FIFO_27[0];
    assign o_Psram_En_To_Sram[28*1 +: 1] = Psram_En_To_Sram_FIFO_28[0];
    assign o_Psram_En_To_Sram[29*1 +: 1] = Psram_En_To_Sram_FIFO_29[0];
    assign o_Psram_En_To_Sram[30*1 +: 1] = Psram_En_To_Sram_FIFO_30[0];
    assign o_Psram_En_To_Sram[31*1 +: 1] = Psram_En_To_Sram_FIFO_31[0];

    // Psram_Valid_To_Systolic Assignments
    assign o_Psram_Valid_To_Systolic[0*1 +: 1] = i_Psram_Valid_1buf;
    assign o_Psram_Valid_To_Systolic[1*1 +: 1] = Psram_Valid_To_Systolic_FIFO_1[0];
    assign o_Psram_Valid_To_Systolic[2*1 +: 1] = Psram_Valid_To_Systolic_FIFO_2[0];
    assign o_Psram_Valid_To_Systolic[3*1 +: 1] = Psram_Valid_To_Systolic_FIFO_3[0];
    assign o_Psram_Valid_To_Systolic[4*1 +: 1] = Psram_Valid_To_Systolic_FIFO_4[0];
    assign o_Psram_Valid_To_Systolic[5*1 +: 1] = Psram_Valid_To_Systolic_FIFO_5[0];
    assign o_Psram_Valid_To_Systolic[6*1 +: 1] = Psram_Valid_To_Systolic_FIFO_6[0];
    assign o_Psram_Valid_To_Systolic[7*1 +: 1] = Psram_Valid_To_Systolic_FIFO_7[0];
    assign o_Psram_Valid_To_Systolic[8*1 +: 1] = Psram_Valid_To_Systolic_FIFO_8[0];
    assign o_Psram_Valid_To_Systolic[9*1 +: 1] = Psram_Valid_To_Systolic_FIFO_9[0];
    assign o_Psram_Valid_To_Systolic[10*1 +: 1] = Psram_Valid_To_Systolic_FIFO_10[0];
    assign o_Psram_Valid_To_Systolic[11*1 +: 1] = Psram_Valid_To_Systolic_FIFO_11[0];
    assign o_Psram_Valid_To_Systolic[12*1 +: 1] = Psram_Valid_To_Systolic_FIFO_12[0];
    assign o_Psram_Valid_To_Systolic[13*1 +: 1] = Psram_Valid_To_Systolic_FIFO_13[0];
    assign o_Psram_Valid_To_Systolic[14*1 +: 1] = Psram_Valid_To_Systolic_FIFO_14[0];
    assign o_Psram_Valid_To_Systolic[15*1 +: 1] = Psram_Valid_To_Systolic_FIFO_15[0];
    assign o_Psram_Valid_To_Systolic[16*1 +: 1] = Psram_Valid_To_Systolic_FIFO_16[0];
    assign o_Psram_Valid_To_Systolic[17*1 +: 1] = Psram_Valid_To_Systolic_FIFO_17[0];
    assign o_Psram_Valid_To_Systolic[18*1 +: 1] = Psram_Valid_To_Systolic_FIFO_18[0];
    assign o_Psram_Valid_To_Systolic[19*1 +: 1] = Psram_Valid_To_Systolic_FIFO_19[0];
    assign o_Psram_Valid_To_Systolic[20*1 +: 1] = Psram_Valid_To_Systolic_FIFO_20[0];
    assign o_Psram_Valid_To_Systolic[21*1 +: 1] = Psram_Valid_To_Systolic_FIFO_21[0];
    assign o_Psram_Valid_To_Systolic[22*1 +: 1] = Psram_Valid_To_Systolic_FIFO_22[0];
    assign o_Psram_Valid_To_Systolic[23*1 +: 1] = Psram_Valid_To_Systolic_FIFO_23[0];
    assign o_Psram_Valid_To_Systolic[24*1 +: 1] = Psram_Valid_To_Systolic_FIFO_24[0];
    assign o_Psram_Valid_To_Systolic[25*1 +: 1] = Psram_Valid_To_Systolic_FIFO_25[0];
    assign o_Psram_Valid_To_Systolic[26*1 +: 1] = Psram_Valid_To_Systolic_FIFO_26[0];
    assign o_Psram_Valid_To_Systolic[27*1 +: 1] = Psram_Valid_To_Systolic_FIFO_27[0];
    assign o_Psram_Valid_To_Systolic[28*1 +: 1] = Psram_Valid_To_Systolic_FIFO_28[0];
    assign o_Psram_Valid_To_Systolic[29*1 +: 1] = Psram_Valid_To_Systolic_FIFO_29[0];
    assign o_Psram_Valid_To_Systolic[30*1 +: 1] = Psram_Valid_To_Systolic_FIFO_30[0];
    assign o_Psram_Valid_To_Systolic[31*1 +: 1] = Psram_Valid_To_Systolic_FIFO_31[0];

    // Psram_Addr_To_Sram Logic
    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_1[0] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_2[0] <= Psram_Addr_To_Sram_FIFO_2[1];
        Psram_Addr_To_Sram_FIFO_3[0] <= Psram_Addr_To_Sram_FIFO_3[1];
        Psram_Addr_To_Sram_FIFO_4[0] <= Psram_Addr_To_Sram_FIFO_4[1];
        Psram_Addr_To_Sram_FIFO_5[0] <= Psram_Addr_To_Sram_FIFO_5[1];
        Psram_Addr_To_Sram_FIFO_6[0] <= Psram_Addr_To_Sram_FIFO_6[1];
        Psram_Addr_To_Sram_FIFO_7[0] <= Psram_Addr_To_Sram_FIFO_7[1];
        Psram_Addr_To_Sram_FIFO_8[0] <= Psram_Addr_To_Sram_FIFO_8[1];
        Psram_Addr_To_Sram_FIFO_9[0] <= Psram_Addr_To_Sram_FIFO_9[1];
        Psram_Addr_To_Sram_FIFO_10[0] <= Psram_Addr_To_Sram_FIFO_10[1];
        Psram_Addr_To_Sram_FIFO_11[0] <= Psram_Addr_To_Sram_FIFO_11[1];
        Psram_Addr_To_Sram_FIFO_12[0] <= Psram_Addr_To_Sram_FIFO_12[1];
        Psram_Addr_To_Sram_FIFO_13[0] <= Psram_Addr_To_Sram_FIFO_13[1];
        Psram_Addr_To_Sram_FIFO_14[0] <= Psram_Addr_To_Sram_FIFO_14[1];
        Psram_Addr_To_Sram_FIFO_15[0] <= Psram_Addr_To_Sram_FIFO_15[1];
        Psram_Addr_To_Sram_FIFO_16[0] <= Psram_Addr_To_Sram_FIFO_16[1];
        Psram_Addr_To_Sram_FIFO_17[0] <= Psram_Addr_To_Sram_FIFO_17[1];
        Psram_Addr_To_Sram_FIFO_18[0] <= Psram_Addr_To_Sram_FIFO_18[1];
        Psram_Addr_To_Sram_FIFO_19[0] <= Psram_Addr_To_Sram_FIFO_19[1];
        Psram_Addr_To_Sram_FIFO_20[0] <= Psram_Addr_To_Sram_FIFO_20[1];
        Psram_Addr_To_Sram_FIFO_21[0] <= Psram_Addr_To_Sram_FIFO_21[1];
        Psram_Addr_To_Sram_FIFO_22[0] <= Psram_Addr_To_Sram_FIFO_22[1];
        Psram_Addr_To_Sram_FIFO_23[0] <= Psram_Addr_To_Sram_FIFO_23[1];
        Psram_Addr_To_Sram_FIFO_24[0] <= Psram_Addr_To_Sram_FIFO_24[1];
        Psram_Addr_To_Sram_FIFO_25[0] <= Psram_Addr_To_Sram_FIFO_25[1];
        Psram_Addr_To_Sram_FIFO_26[0] <= Psram_Addr_To_Sram_FIFO_26[1];
        Psram_Addr_To_Sram_FIFO_27[0] <= Psram_Addr_To_Sram_FIFO_27[1];
        Psram_Addr_To_Sram_FIFO_28[0] <= Psram_Addr_To_Sram_FIFO_28[1];
        Psram_Addr_To_Sram_FIFO_29[0] <= Psram_Addr_To_Sram_FIFO_29[1];
        Psram_Addr_To_Sram_FIFO_30[0] <= Psram_Addr_To_Sram_FIFO_30[1];
        Psram_Addr_To_Sram_FIFO_31[0] <= Psram_Addr_To_Sram_FIFO_31[1];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_2[1] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_3[1] <= Psram_Addr_To_Sram_FIFO_3[2];
        Psram_Addr_To_Sram_FIFO_4[1] <= Psram_Addr_To_Sram_FIFO_4[2];
        Psram_Addr_To_Sram_FIFO_5[1] <= Psram_Addr_To_Sram_FIFO_5[2];
        Psram_Addr_To_Sram_FIFO_6[1] <= Psram_Addr_To_Sram_FIFO_6[2];
        Psram_Addr_To_Sram_FIFO_7[1] <= Psram_Addr_To_Sram_FIFO_7[2];
        Psram_Addr_To_Sram_FIFO_8[1] <= Psram_Addr_To_Sram_FIFO_8[2];
        Psram_Addr_To_Sram_FIFO_9[1] <= Psram_Addr_To_Sram_FIFO_9[2];
        Psram_Addr_To_Sram_FIFO_10[1] <= Psram_Addr_To_Sram_FIFO_10[2];
        Psram_Addr_To_Sram_FIFO_11[1] <= Psram_Addr_To_Sram_FIFO_11[2];
        Psram_Addr_To_Sram_FIFO_12[1] <= Psram_Addr_To_Sram_FIFO_12[2];
        Psram_Addr_To_Sram_FIFO_13[1] <= Psram_Addr_To_Sram_FIFO_13[2];
        Psram_Addr_To_Sram_FIFO_14[1] <= Psram_Addr_To_Sram_FIFO_14[2];
        Psram_Addr_To_Sram_FIFO_15[1] <= Psram_Addr_To_Sram_FIFO_15[2];
        Psram_Addr_To_Sram_FIFO_16[1] <= Psram_Addr_To_Sram_FIFO_16[2];
        Psram_Addr_To_Sram_FIFO_17[1] <= Psram_Addr_To_Sram_FIFO_17[2];
        Psram_Addr_To_Sram_FIFO_18[1] <= Psram_Addr_To_Sram_FIFO_18[2];
        Psram_Addr_To_Sram_FIFO_19[1] <= Psram_Addr_To_Sram_FIFO_19[2];
        Psram_Addr_To_Sram_FIFO_20[1] <= Psram_Addr_To_Sram_FIFO_20[2];
        Psram_Addr_To_Sram_FIFO_21[1] <= Psram_Addr_To_Sram_FIFO_21[2];
        Psram_Addr_To_Sram_FIFO_22[1] <= Psram_Addr_To_Sram_FIFO_22[2];
        Psram_Addr_To_Sram_FIFO_23[1] <= Psram_Addr_To_Sram_FIFO_23[2];
        Psram_Addr_To_Sram_FIFO_24[1] <= Psram_Addr_To_Sram_FIFO_24[2];
        Psram_Addr_To_Sram_FIFO_25[1] <= Psram_Addr_To_Sram_FIFO_25[2];
        Psram_Addr_To_Sram_FIFO_26[1] <= Psram_Addr_To_Sram_FIFO_26[2];
        Psram_Addr_To_Sram_FIFO_27[1] <= Psram_Addr_To_Sram_FIFO_27[2];
        Psram_Addr_To_Sram_FIFO_28[1] <= Psram_Addr_To_Sram_FIFO_28[2];
        Psram_Addr_To_Sram_FIFO_29[1] <= Psram_Addr_To_Sram_FIFO_29[2];
        Psram_Addr_To_Sram_FIFO_30[1] <= Psram_Addr_To_Sram_FIFO_30[2];
        Psram_Addr_To_Sram_FIFO_31[1] <= Psram_Addr_To_Sram_FIFO_31[2];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_3[2] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_4[2] <= Psram_Addr_To_Sram_FIFO_4[3];
        Psram_Addr_To_Sram_FIFO_5[2] <= Psram_Addr_To_Sram_FIFO_5[3];
        Psram_Addr_To_Sram_FIFO_6[2] <= Psram_Addr_To_Sram_FIFO_6[3];
        Psram_Addr_To_Sram_FIFO_7[2] <= Psram_Addr_To_Sram_FIFO_7[3];
        Psram_Addr_To_Sram_FIFO_8[2] <= Psram_Addr_To_Sram_FIFO_8[3];
        Psram_Addr_To_Sram_FIFO_9[2] <= Psram_Addr_To_Sram_FIFO_9[3];
        Psram_Addr_To_Sram_FIFO_10[2] <= Psram_Addr_To_Sram_FIFO_10[3];
        Psram_Addr_To_Sram_FIFO_11[2] <= Psram_Addr_To_Sram_FIFO_11[3];
        Psram_Addr_To_Sram_FIFO_12[2] <= Psram_Addr_To_Sram_FIFO_12[3];
        Psram_Addr_To_Sram_FIFO_13[2] <= Psram_Addr_To_Sram_FIFO_13[3];
        Psram_Addr_To_Sram_FIFO_14[2] <= Psram_Addr_To_Sram_FIFO_14[3];
        Psram_Addr_To_Sram_FIFO_15[2] <= Psram_Addr_To_Sram_FIFO_15[3];
        Psram_Addr_To_Sram_FIFO_16[2] <= Psram_Addr_To_Sram_FIFO_16[3];
        Psram_Addr_To_Sram_FIFO_17[2] <= Psram_Addr_To_Sram_FIFO_17[3];
        Psram_Addr_To_Sram_FIFO_18[2] <= Psram_Addr_To_Sram_FIFO_18[3];
        Psram_Addr_To_Sram_FIFO_19[2] <= Psram_Addr_To_Sram_FIFO_19[3];
        Psram_Addr_To_Sram_FIFO_20[2] <= Psram_Addr_To_Sram_FIFO_20[3];
        Psram_Addr_To_Sram_FIFO_21[2] <= Psram_Addr_To_Sram_FIFO_21[3];
        Psram_Addr_To_Sram_FIFO_22[2] <= Psram_Addr_To_Sram_FIFO_22[3];
        Psram_Addr_To_Sram_FIFO_23[2] <= Psram_Addr_To_Sram_FIFO_23[3];
        Psram_Addr_To_Sram_FIFO_24[2] <= Psram_Addr_To_Sram_FIFO_24[3];
        Psram_Addr_To_Sram_FIFO_25[2] <= Psram_Addr_To_Sram_FIFO_25[3];
        Psram_Addr_To_Sram_FIFO_26[2] <= Psram_Addr_To_Sram_FIFO_26[3];
        Psram_Addr_To_Sram_FIFO_27[2] <= Psram_Addr_To_Sram_FIFO_27[3];
        Psram_Addr_To_Sram_FIFO_28[2] <= Psram_Addr_To_Sram_FIFO_28[3];
        Psram_Addr_To_Sram_FIFO_29[2] <= Psram_Addr_To_Sram_FIFO_29[3];
        Psram_Addr_To_Sram_FIFO_30[2] <= Psram_Addr_To_Sram_FIFO_30[3];
        Psram_Addr_To_Sram_FIFO_31[2] <= Psram_Addr_To_Sram_FIFO_31[3];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_4[3] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_5[3] <= Psram_Addr_To_Sram_FIFO_5[4];
        Psram_Addr_To_Sram_FIFO_6[3] <= Psram_Addr_To_Sram_FIFO_6[4];
        Psram_Addr_To_Sram_FIFO_7[3] <= Psram_Addr_To_Sram_FIFO_7[4];
        Psram_Addr_To_Sram_FIFO_8[3] <= Psram_Addr_To_Sram_FIFO_8[4];
        Psram_Addr_To_Sram_FIFO_9[3] <= Psram_Addr_To_Sram_FIFO_9[4];
        Psram_Addr_To_Sram_FIFO_10[3] <= Psram_Addr_To_Sram_FIFO_10[4];
        Psram_Addr_To_Sram_FIFO_11[3] <= Psram_Addr_To_Sram_FIFO_11[4];
        Psram_Addr_To_Sram_FIFO_12[3] <= Psram_Addr_To_Sram_FIFO_12[4];
        Psram_Addr_To_Sram_FIFO_13[3] <= Psram_Addr_To_Sram_FIFO_13[4];
        Psram_Addr_To_Sram_FIFO_14[3] <= Psram_Addr_To_Sram_FIFO_14[4];
        Psram_Addr_To_Sram_FIFO_15[3] <= Psram_Addr_To_Sram_FIFO_15[4];
        Psram_Addr_To_Sram_FIFO_16[3] <= Psram_Addr_To_Sram_FIFO_16[4];
        Psram_Addr_To_Sram_FIFO_17[3] <= Psram_Addr_To_Sram_FIFO_17[4];
        Psram_Addr_To_Sram_FIFO_18[3] <= Psram_Addr_To_Sram_FIFO_18[4];
        Psram_Addr_To_Sram_FIFO_19[3] <= Psram_Addr_To_Sram_FIFO_19[4];
        Psram_Addr_To_Sram_FIFO_20[3] <= Psram_Addr_To_Sram_FIFO_20[4];
        Psram_Addr_To_Sram_FIFO_21[3] <= Psram_Addr_To_Sram_FIFO_21[4];
        Psram_Addr_To_Sram_FIFO_22[3] <= Psram_Addr_To_Sram_FIFO_22[4];
        Psram_Addr_To_Sram_FIFO_23[3] <= Psram_Addr_To_Sram_FIFO_23[4];
        Psram_Addr_To_Sram_FIFO_24[3] <= Psram_Addr_To_Sram_FIFO_24[4];
        Psram_Addr_To_Sram_FIFO_25[3] <= Psram_Addr_To_Sram_FIFO_25[4];
        Psram_Addr_To_Sram_FIFO_26[3] <= Psram_Addr_To_Sram_FIFO_26[4];
        Psram_Addr_To_Sram_FIFO_27[3] <= Psram_Addr_To_Sram_FIFO_27[4];
        Psram_Addr_To_Sram_FIFO_28[3] <= Psram_Addr_To_Sram_FIFO_28[4];
        Psram_Addr_To_Sram_FIFO_29[3] <= Psram_Addr_To_Sram_FIFO_29[4];
        Psram_Addr_To_Sram_FIFO_30[3] <= Psram_Addr_To_Sram_FIFO_30[4];
        Psram_Addr_To_Sram_FIFO_31[3] <= Psram_Addr_To_Sram_FIFO_31[4];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_5[4] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_6[4] <= Psram_Addr_To_Sram_FIFO_6[5];
        Psram_Addr_To_Sram_FIFO_7[4] <= Psram_Addr_To_Sram_FIFO_7[5];
        Psram_Addr_To_Sram_FIFO_8[4] <= Psram_Addr_To_Sram_FIFO_8[5];
        Psram_Addr_To_Sram_FIFO_9[4] <= Psram_Addr_To_Sram_FIFO_9[5];
        Psram_Addr_To_Sram_FIFO_10[4] <= Psram_Addr_To_Sram_FIFO_10[5];
        Psram_Addr_To_Sram_FIFO_11[4] <= Psram_Addr_To_Sram_FIFO_11[5];
        Psram_Addr_To_Sram_FIFO_12[4] <= Psram_Addr_To_Sram_FIFO_12[5];
        Psram_Addr_To_Sram_FIFO_13[4] <= Psram_Addr_To_Sram_FIFO_13[5];
        Psram_Addr_To_Sram_FIFO_14[4] <= Psram_Addr_To_Sram_FIFO_14[5];
        Psram_Addr_To_Sram_FIFO_15[4] <= Psram_Addr_To_Sram_FIFO_15[5];
        Psram_Addr_To_Sram_FIFO_16[4] <= Psram_Addr_To_Sram_FIFO_16[5];
        Psram_Addr_To_Sram_FIFO_17[4] <= Psram_Addr_To_Sram_FIFO_17[5];
        Psram_Addr_To_Sram_FIFO_18[4] <= Psram_Addr_To_Sram_FIFO_18[5];
        Psram_Addr_To_Sram_FIFO_19[4] <= Psram_Addr_To_Sram_FIFO_19[5];
        Psram_Addr_To_Sram_FIFO_20[4] <= Psram_Addr_To_Sram_FIFO_20[5];
        Psram_Addr_To_Sram_FIFO_21[4] <= Psram_Addr_To_Sram_FIFO_21[5];
        Psram_Addr_To_Sram_FIFO_22[4] <= Psram_Addr_To_Sram_FIFO_22[5];
        Psram_Addr_To_Sram_FIFO_23[4] <= Psram_Addr_To_Sram_FIFO_23[5];
        Psram_Addr_To_Sram_FIFO_24[4] <= Psram_Addr_To_Sram_FIFO_24[5];
        Psram_Addr_To_Sram_FIFO_25[4] <= Psram_Addr_To_Sram_FIFO_25[5];
        Psram_Addr_To_Sram_FIFO_26[4] <= Psram_Addr_To_Sram_FIFO_26[5];
        Psram_Addr_To_Sram_FIFO_27[4] <= Psram_Addr_To_Sram_FIFO_27[5];
        Psram_Addr_To_Sram_FIFO_28[4] <= Psram_Addr_To_Sram_FIFO_28[5];
        Psram_Addr_To_Sram_FIFO_29[4] <= Psram_Addr_To_Sram_FIFO_29[5];
        Psram_Addr_To_Sram_FIFO_30[4] <= Psram_Addr_To_Sram_FIFO_30[5];
        Psram_Addr_To_Sram_FIFO_31[4] <= Psram_Addr_To_Sram_FIFO_31[5];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_6[5] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_7[5] <= Psram_Addr_To_Sram_FIFO_7[6];
        Psram_Addr_To_Sram_FIFO_8[5] <= Psram_Addr_To_Sram_FIFO_8[6];
        Psram_Addr_To_Sram_FIFO_9[5] <= Psram_Addr_To_Sram_FIFO_9[6];
        Psram_Addr_To_Sram_FIFO_10[5] <= Psram_Addr_To_Sram_FIFO_10[6];
        Psram_Addr_To_Sram_FIFO_11[5] <= Psram_Addr_To_Sram_FIFO_11[6];
        Psram_Addr_To_Sram_FIFO_12[5] <= Psram_Addr_To_Sram_FIFO_12[6];
        Psram_Addr_To_Sram_FIFO_13[5] <= Psram_Addr_To_Sram_FIFO_13[6];
        Psram_Addr_To_Sram_FIFO_14[5] <= Psram_Addr_To_Sram_FIFO_14[6];
        Psram_Addr_To_Sram_FIFO_15[5] <= Psram_Addr_To_Sram_FIFO_15[6];
        Psram_Addr_To_Sram_FIFO_16[5] <= Psram_Addr_To_Sram_FIFO_16[6];
        Psram_Addr_To_Sram_FIFO_17[5] <= Psram_Addr_To_Sram_FIFO_17[6];
        Psram_Addr_To_Sram_FIFO_18[5] <= Psram_Addr_To_Sram_FIFO_18[6];
        Psram_Addr_To_Sram_FIFO_19[5] <= Psram_Addr_To_Sram_FIFO_19[6];
        Psram_Addr_To_Sram_FIFO_20[5] <= Psram_Addr_To_Sram_FIFO_20[6];
        Psram_Addr_To_Sram_FIFO_21[5] <= Psram_Addr_To_Sram_FIFO_21[6];
        Psram_Addr_To_Sram_FIFO_22[5] <= Psram_Addr_To_Sram_FIFO_22[6];
        Psram_Addr_To_Sram_FIFO_23[5] <= Psram_Addr_To_Sram_FIFO_23[6];
        Psram_Addr_To_Sram_FIFO_24[5] <= Psram_Addr_To_Sram_FIFO_24[6];
        Psram_Addr_To_Sram_FIFO_25[5] <= Psram_Addr_To_Sram_FIFO_25[6];
        Psram_Addr_To_Sram_FIFO_26[5] <= Psram_Addr_To_Sram_FIFO_26[6];
        Psram_Addr_To_Sram_FIFO_27[5] <= Psram_Addr_To_Sram_FIFO_27[6];
        Psram_Addr_To_Sram_FIFO_28[5] <= Psram_Addr_To_Sram_FIFO_28[6];
        Psram_Addr_To_Sram_FIFO_29[5] <= Psram_Addr_To_Sram_FIFO_29[6];
        Psram_Addr_To_Sram_FIFO_30[5] <= Psram_Addr_To_Sram_FIFO_30[6];
        Psram_Addr_To_Sram_FIFO_31[5] <= Psram_Addr_To_Sram_FIFO_31[6];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_7[6] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_8[6] <= Psram_Addr_To_Sram_FIFO_8[7];
        Psram_Addr_To_Sram_FIFO_9[6] <= Psram_Addr_To_Sram_FIFO_9[7];
        Psram_Addr_To_Sram_FIFO_10[6] <= Psram_Addr_To_Sram_FIFO_10[7];
        Psram_Addr_To_Sram_FIFO_11[6] <= Psram_Addr_To_Sram_FIFO_11[7];
        Psram_Addr_To_Sram_FIFO_12[6] <= Psram_Addr_To_Sram_FIFO_12[7];
        Psram_Addr_To_Sram_FIFO_13[6] <= Psram_Addr_To_Sram_FIFO_13[7];
        Psram_Addr_To_Sram_FIFO_14[6] <= Psram_Addr_To_Sram_FIFO_14[7];
        Psram_Addr_To_Sram_FIFO_15[6] <= Psram_Addr_To_Sram_FIFO_15[7];
        Psram_Addr_To_Sram_FIFO_16[6] <= Psram_Addr_To_Sram_FIFO_16[7];
        Psram_Addr_To_Sram_FIFO_17[6] <= Psram_Addr_To_Sram_FIFO_17[7];
        Psram_Addr_To_Sram_FIFO_18[6] <= Psram_Addr_To_Sram_FIFO_18[7];
        Psram_Addr_To_Sram_FIFO_19[6] <= Psram_Addr_To_Sram_FIFO_19[7];
        Psram_Addr_To_Sram_FIFO_20[6] <= Psram_Addr_To_Sram_FIFO_20[7];
        Psram_Addr_To_Sram_FIFO_21[6] <= Psram_Addr_To_Sram_FIFO_21[7];
        Psram_Addr_To_Sram_FIFO_22[6] <= Psram_Addr_To_Sram_FIFO_22[7];
        Psram_Addr_To_Sram_FIFO_23[6] <= Psram_Addr_To_Sram_FIFO_23[7];
        Psram_Addr_To_Sram_FIFO_24[6] <= Psram_Addr_To_Sram_FIFO_24[7];
        Psram_Addr_To_Sram_FIFO_25[6] <= Psram_Addr_To_Sram_FIFO_25[7];
        Psram_Addr_To_Sram_FIFO_26[6] <= Psram_Addr_To_Sram_FIFO_26[7];
        Psram_Addr_To_Sram_FIFO_27[6] <= Psram_Addr_To_Sram_FIFO_27[7];
        Psram_Addr_To_Sram_FIFO_28[6] <= Psram_Addr_To_Sram_FIFO_28[7];
        Psram_Addr_To_Sram_FIFO_29[6] <= Psram_Addr_To_Sram_FIFO_29[7];
        Psram_Addr_To_Sram_FIFO_30[6] <= Psram_Addr_To_Sram_FIFO_30[7];
        Psram_Addr_To_Sram_FIFO_31[6] <= Psram_Addr_To_Sram_FIFO_31[7];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_8[7] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_9[7] <= Psram_Addr_To_Sram_FIFO_9[8];
        Psram_Addr_To_Sram_FIFO_10[7] <= Psram_Addr_To_Sram_FIFO_10[8];
        Psram_Addr_To_Sram_FIFO_11[7] <= Psram_Addr_To_Sram_FIFO_11[8];
        Psram_Addr_To_Sram_FIFO_12[7] <= Psram_Addr_To_Sram_FIFO_12[8];
        Psram_Addr_To_Sram_FIFO_13[7] <= Psram_Addr_To_Sram_FIFO_13[8];
        Psram_Addr_To_Sram_FIFO_14[7] <= Psram_Addr_To_Sram_FIFO_14[8];
        Psram_Addr_To_Sram_FIFO_15[7] <= Psram_Addr_To_Sram_FIFO_15[8];
        Psram_Addr_To_Sram_FIFO_16[7] <= Psram_Addr_To_Sram_FIFO_16[8];
        Psram_Addr_To_Sram_FIFO_17[7] <= Psram_Addr_To_Sram_FIFO_17[8];
        Psram_Addr_To_Sram_FIFO_18[7] <= Psram_Addr_To_Sram_FIFO_18[8];
        Psram_Addr_To_Sram_FIFO_19[7] <= Psram_Addr_To_Sram_FIFO_19[8];
        Psram_Addr_To_Sram_FIFO_20[7] <= Psram_Addr_To_Sram_FIFO_20[8];
        Psram_Addr_To_Sram_FIFO_21[7] <= Psram_Addr_To_Sram_FIFO_21[8];
        Psram_Addr_To_Sram_FIFO_22[7] <= Psram_Addr_To_Sram_FIFO_22[8];
        Psram_Addr_To_Sram_FIFO_23[7] <= Psram_Addr_To_Sram_FIFO_23[8];
        Psram_Addr_To_Sram_FIFO_24[7] <= Psram_Addr_To_Sram_FIFO_24[8];
        Psram_Addr_To_Sram_FIFO_25[7] <= Psram_Addr_To_Sram_FIFO_25[8];
        Psram_Addr_To_Sram_FIFO_26[7] <= Psram_Addr_To_Sram_FIFO_26[8];
        Psram_Addr_To_Sram_FIFO_27[7] <= Psram_Addr_To_Sram_FIFO_27[8];
        Psram_Addr_To_Sram_FIFO_28[7] <= Psram_Addr_To_Sram_FIFO_28[8];
        Psram_Addr_To_Sram_FIFO_29[7] <= Psram_Addr_To_Sram_FIFO_29[8];
        Psram_Addr_To_Sram_FIFO_30[7] <= Psram_Addr_To_Sram_FIFO_30[8];
        Psram_Addr_To_Sram_FIFO_31[7] <= Psram_Addr_To_Sram_FIFO_31[8];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_9[8] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_10[8] <= Psram_Addr_To_Sram_FIFO_10[9];
        Psram_Addr_To_Sram_FIFO_11[8] <= Psram_Addr_To_Sram_FIFO_11[9];
        Psram_Addr_To_Sram_FIFO_12[8] <= Psram_Addr_To_Sram_FIFO_12[9];
        Psram_Addr_To_Sram_FIFO_13[8] <= Psram_Addr_To_Sram_FIFO_13[9];
        Psram_Addr_To_Sram_FIFO_14[8] <= Psram_Addr_To_Sram_FIFO_14[9];
        Psram_Addr_To_Sram_FIFO_15[8] <= Psram_Addr_To_Sram_FIFO_15[9];
        Psram_Addr_To_Sram_FIFO_16[8] <= Psram_Addr_To_Sram_FIFO_16[9];
        Psram_Addr_To_Sram_FIFO_17[8] <= Psram_Addr_To_Sram_FIFO_17[9];
        Psram_Addr_To_Sram_FIFO_18[8] <= Psram_Addr_To_Sram_FIFO_18[9];
        Psram_Addr_To_Sram_FIFO_19[8] <= Psram_Addr_To_Sram_FIFO_19[9];
        Psram_Addr_To_Sram_FIFO_20[8] <= Psram_Addr_To_Sram_FIFO_20[9];
        Psram_Addr_To_Sram_FIFO_21[8] <= Psram_Addr_To_Sram_FIFO_21[9];
        Psram_Addr_To_Sram_FIFO_22[8] <= Psram_Addr_To_Sram_FIFO_22[9];
        Psram_Addr_To_Sram_FIFO_23[8] <= Psram_Addr_To_Sram_FIFO_23[9];
        Psram_Addr_To_Sram_FIFO_24[8] <= Psram_Addr_To_Sram_FIFO_24[9];
        Psram_Addr_To_Sram_FIFO_25[8] <= Psram_Addr_To_Sram_FIFO_25[9];
        Psram_Addr_To_Sram_FIFO_26[8] <= Psram_Addr_To_Sram_FIFO_26[9];
        Psram_Addr_To_Sram_FIFO_27[8] <= Psram_Addr_To_Sram_FIFO_27[9];
        Psram_Addr_To_Sram_FIFO_28[8] <= Psram_Addr_To_Sram_FIFO_28[9];
        Psram_Addr_To_Sram_FIFO_29[8] <= Psram_Addr_To_Sram_FIFO_29[9];
        Psram_Addr_To_Sram_FIFO_30[8] <= Psram_Addr_To_Sram_FIFO_30[9];
        Psram_Addr_To_Sram_FIFO_31[8] <= Psram_Addr_To_Sram_FIFO_31[9];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_10[9] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_11[9] <= Psram_Addr_To_Sram_FIFO_11[10];
        Psram_Addr_To_Sram_FIFO_12[9] <= Psram_Addr_To_Sram_FIFO_12[10];
        Psram_Addr_To_Sram_FIFO_13[9] <= Psram_Addr_To_Sram_FIFO_13[10];
        Psram_Addr_To_Sram_FIFO_14[9] <= Psram_Addr_To_Sram_FIFO_14[10];
        Psram_Addr_To_Sram_FIFO_15[9] <= Psram_Addr_To_Sram_FIFO_15[10];
        Psram_Addr_To_Sram_FIFO_16[9] <= Psram_Addr_To_Sram_FIFO_16[10];
        Psram_Addr_To_Sram_FIFO_17[9] <= Psram_Addr_To_Sram_FIFO_17[10];
        Psram_Addr_To_Sram_FIFO_18[9] <= Psram_Addr_To_Sram_FIFO_18[10];
        Psram_Addr_To_Sram_FIFO_19[9] <= Psram_Addr_To_Sram_FIFO_19[10];
        Psram_Addr_To_Sram_FIFO_20[9] <= Psram_Addr_To_Sram_FIFO_20[10];
        Psram_Addr_To_Sram_FIFO_21[9] <= Psram_Addr_To_Sram_FIFO_21[10];
        Psram_Addr_To_Sram_FIFO_22[9] <= Psram_Addr_To_Sram_FIFO_22[10];
        Psram_Addr_To_Sram_FIFO_23[9] <= Psram_Addr_To_Sram_FIFO_23[10];
        Psram_Addr_To_Sram_FIFO_24[9] <= Psram_Addr_To_Sram_FIFO_24[10];
        Psram_Addr_To_Sram_FIFO_25[9] <= Psram_Addr_To_Sram_FIFO_25[10];
        Psram_Addr_To_Sram_FIFO_26[9] <= Psram_Addr_To_Sram_FIFO_26[10];
        Psram_Addr_To_Sram_FIFO_27[9] <= Psram_Addr_To_Sram_FIFO_27[10];
        Psram_Addr_To_Sram_FIFO_28[9] <= Psram_Addr_To_Sram_FIFO_28[10];
        Psram_Addr_To_Sram_FIFO_29[9] <= Psram_Addr_To_Sram_FIFO_29[10];
        Psram_Addr_To_Sram_FIFO_30[9] <= Psram_Addr_To_Sram_FIFO_30[10];
        Psram_Addr_To_Sram_FIFO_31[9] <= Psram_Addr_To_Sram_FIFO_31[10];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_11[10] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_12[10] <= Psram_Addr_To_Sram_FIFO_12[11];
        Psram_Addr_To_Sram_FIFO_13[10] <= Psram_Addr_To_Sram_FIFO_13[11];
        Psram_Addr_To_Sram_FIFO_14[10] <= Psram_Addr_To_Sram_FIFO_14[11];
        Psram_Addr_To_Sram_FIFO_15[10] <= Psram_Addr_To_Sram_FIFO_15[11];
        Psram_Addr_To_Sram_FIFO_16[10] <= Psram_Addr_To_Sram_FIFO_16[11];
        Psram_Addr_To_Sram_FIFO_17[10] <= Psram_Addr_To_Sram_FIFO_17[11];
        Psram_Addr_To_Sram_FIFO_18[10] <= Psram_Addr_To_Sram_FIFO_18[11];
        Psram_Addr_To_Sram_FIFO_19[10] <= Psram_Addr_To_Sram_FIFO_19[11];
        Psram_Addr_To_Sram_FIFO_20[10] <= Psram_Addr_To_Sram_FIFO_20[11];
        Psram_Addr_To_Sram_FIFO_21[10] <= Psram_Addr_To_Sram_FIFO_21[11];
        Psram_Addr_To_Sram_FIFO_22[10] <= Psram_Addr_To_Sram_FIFO_22[11];
        Psram_Addr_To_Sram_FIFO_23[10] <= Psram_Addr_To_Sram_FIFO_23[11];
        Psram_Addr_To_Sram_FIFO_24[10] <= Psram_Addr_To_Sram_FIFO_24[11];
        Psram_Addr_To_Sram_FIFO_25[10] <= Psram_Addr_To_Sram_FIFO_25[11];
        Psram_Addr_To_Sram_FIFO_26[10] <= Psram_Addr_To_Sram_FIFO_26[11];
        Psram_Addr_To_Sram_FIFO_27[10] <= Psram_Addr_To_Sram_FIFO_27[11];
        Psram_Addr_To_Sram_FIFO_28[10] <= Psram_Addr_To_Sram_FIFO_28[11];
        Psram_Addr_To_Sram_FIFO_29[10] <= Psram_Addr_To_Sram_FIFO_29[11];
        Psram_Addr_To_Sram_FIFO_30[10] <= Psram_Addr_To_Sram_FIFO_30[11];
        Psram_Addr_To_Sram_FIFO_31[10] <= Psram_Addr_To_Sram_FIFO_31[11];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_12[11] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_13[11] <= Psram_Addr_To_Sram_FIFO_13[12];
        Psram_Addr_To_Sram_FIFO_14[11] <= Psram_Addr_To_Sram_FIFO_14[12];
        Psram_Addr_To_Sram_FIFO_15[11] <= Psram_Addr_To_Sram_FIFO_15[12];
        Psram_Addr_To_Sram_FIFO_16[11] <= Psram_Addr_To_Sram_FIFO_16[12];
        Psram_Addr_To_Sram_FIFO_17[11] <= Psram_Addr_To_Sram_FIFO_17[12];
        Psram_Addr_To_Sram_FIFO_18[11] <= Psram_Addr_To_Sram_FIFO_18[12];
        Psram_Addr_To_Sram_FIFO_19[11] <= Psram_Addr_To_Sram_FIFO_19[12];
        Psram_Addr_To_Sram_FIFO_20[11] <= Psram_Addr_To_Sram_FIFO_20[12];
        Psram_Addr_To_Sram_FIFO_21[11] <= Psram_Addr_To_Sram_FIFO_21[12];
        Psram_Addr_To_Sram_FIFO_22[11] <= Psram_Addr_To_Sram_FIFO_22[12];
        Psram_Addr_To_Sram_FIFO_23[11] <= Psram_Addr_To_Sram_FIFO_23[12];
        Psram_Addr_To_Sram_FIFO_24[11] <= Psram_Addr_To_Sram_FIFO_24[12];
        Psram_Addr_To_Sram_FIFO_25[11] <= Psram_Addr_To_Sram_FIFO_25[12];
        Psram_Addr_To_Sram_FIFO_26[11] <= Psram_Addr_To_Sram_FIFO_26[12];
        Psram_Addr_To_Sram_FIFO_27[11] <= Psram_Addr_To_Sram_FIFO_27[12];
        Psram_Addr_To_Sram_FIFO_28[11] <= Psram_Addr_To_Sram_FIFO_28[12];
        Psram_Addr_To_Sram_FIFO_29[11] <= Psram_Addr_To_Sram_FIFO_29[12];
        Psram_Addr_To_Sram_FIFO_30[11] <= Psram_Addr_To_Sram_FIFO_30[12];
        Psram_Addr_To_Sram_FIFO_31[11] <= Psram_Addr_To_Sram_FIFO_31[12];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_13[12] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_14[12] <= Psram_Addr_To_Sram_FIFO_14[13];
        Psram_Addr_To_Sram_FIFO_15[12] <= Psram_Addr_To_Sram_FIFO_15[13];
        Psram_Addr_To_Sram_FIFO_16[12] <= Psram_Addr_To_Sram_FIFO_16[13];
        Psram_Addr_To_Sram_FIFO_17[12] <= Psram_Addr_To_Sram_FIFO_17[13];
        Psram_Addr_To_Sram_FIFO_18[12] <= Psram_Addr_To_Sram_FIFO_18[13];
        Psram_Addr_To_Sram_FIFO_19[12] <= Psram_Addr_To_Sram_FIFO_19[13];
        Psram_Addr_To_Sram_FIFO_20[12] <= Psram_Addr_To_Sram_FIFO_20[13];
        Psram_Addr_To_Sram_FIFO_21[12] <= Psram_Addr_To_Sram_FIFO_21[13];
        Psram_Addr_To_Sram_FIFO_22[12] <= Psram_Addr_To_Sram_FIFO_22[13];
        Psram_Addr_To_Sram_FIFO_23[12] <= Psram_Addr_To_Sram_FIFO_23[13];
        Psram_Addr_To_Sram_FIFO_24[12] <= Psram_Addr_To_Sram_FIFO_24[13];
        Psram_Addr_To_Sram_FIFO_25[12] <= Psram_Addr_To_Sram_FIFO_25[13];
        Psram_Addr_To_Sram_FIFO_26[12] <= Psram_Addr_To_Sram_FIFO_26[13];
        Psram_Addr_To_Sram_FIFO_27[12] <= Psram_Addr_To_Sram_FIFO_27[13];
        Psram_Addr_To_Sram_FIFO_28[12] <= Psram_Addr_To_Sram_FIFO_28[13];
        Psram_Addr_To_Sram_FIFO_29[12] <= Psram_Addr_To_Sram_FIFO_29[13];
        Psram_Addr_To_Sram_FIFO_30[12] <= Psram_Addr_To_Sram_FIFO_30[13];
        Psram_Addr_To_Sram_FIFO_31[12] <= Psram_Addr_To_Sram_FIFO_31[13];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_14[13] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_15[13] <= Psram_Addr_To_Sram_FIFO_15[14];
        Psram_Addr_To_Sram_FIFO_16[13] <= Psram_Addr_To_Sram_FIFO_16[14];
        Psram_Addr_To_Sram_FIFO_17[13] <= Psram_Addr_To_Sram_FIFO_17[14];
        Psram_Addr_To_Sram_FIFO_18[13] <= Psram_Addr_To_Sram_FIFO_18[14];
        Psram_Addr_To_Sram_FIFO_19[13] <= Psram_Addr_To_Sram_FIFO_19[14];
        Psram_Addr_To_Sram_FIFO_20[13] <= Psram_Addr_To_Sram_FIFO_20[14];
        Psram_Addr_To_Sram_FIFO_21[13] <= Psram_Addr_To_Sram_FIFO_21[14];
        Psram_Addr_To_Sram_FIFO_22[13] <= Psram_Addr_To_Sram_FIFO_22[14];
        Psram_Addr_To_Sram_FIFO_23[13] <= Psram_Addr_To_Sram_FIFO_23[14];
        Psram_Addr_To_Sram_FIFO_24[13] <= Psram_Addr_To_Sram_FIFO_24[14];
        Psram_Addr_To_Sram_FIFO_25[13] <= Psram_Addr_To_Sram_FIFO_25[14];
        Psram_Addr_To_Sram_FIFO_26[13] <= Psram_Addr_To_Sram_FIFO_26[14];
        Psram_Addr_To_Sram_FIFO_27[13] <= Psram_Addr_To_Sram_FIFO_27[14];
        Psram_Addr_To_Sram_FIFO_28[13] <= Psram_Addr_To_Sram_FIFO_28[14];
        Psram_Addr_To_Sram_FIFO_29[13] <= Psram_Addr_To_Sram_FIFO_29[14];
        Psram_Addr_To_Sram_FIFO_30[13] <= Psram_Addr_To_Sram_FIFO_30[14];
        Psram_Addr_To_Sram_FIFO_31[13] <= Psram_Addr_To_Sram_FIFO_31[14];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_15[14] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_16[14] <= Psram_Addr_To_Sram_FIFO_16[15];
        Psram_Addr_To_Sram_FIFO_17[14] <= Psram_Addr_To_Sram_FIFO_17[15];
        Psram_Addr_To_Sram_FIFO_18[14] <= Psram_Addr_To_Sram_FIFO_18[15];
        Psram_Addr_To_Sram_FIFO_19[14] <= Psram_Addr_To_Sram_FIFO_19[15];
        Psram_Addr_To_Sram_FIFO_20[14] <= Psram_Addr_To_Sram_FIFO_20[15];
        Psram_Addr_To_Sram_FIFO_21[14] <= Psram_Addr_To_Sram_FIFO_21[15];
        Psram_Addr_To_Sram_FIFO_22[14] <= Psram_Addr_To_Sram_FIFO_22[15];
        Psram_Addr_To_Sram_FIFO_23[14] <= Psram_Addr_To_Sram_FIFO_23[15];
        Psram_Addr_To_Sram_FIFO_24[14] <= Psram_Addr_To_Sram_FIFO_24[15];
        Psram_Addr_To_Sram_FIFO_25[14] <= Psram_Addr_To_Sram_FIFO_25[15];
        Psram_Addr_To_Sram_FIFO_26[14] <= Psram_Addr_To_Sram_FIFO_26[15];
        Psram_Addr_To_Sram_FIFO_27[14] <= Psram_Addr_To_Sram_FIFO_27[15];
        Psram_Addr_To_Sram_FIFO_28[14] <= Psram_Addr_To_Sram_FIFO_28[15];
        Psram_Addr_To_Sram_FIFO_29[14] <= Psram_Addr_To_Sram_FIFO_29[15];
        Psram_Addr_To_Sram_FIFO_30[14] <= Psram_Addr_To_Sram_FIFO_30[15];
        Psram_Addr_To_Sram_FIFO_31[14] <= Psram_Addr_To_Sram_FIFO_31[15];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_16[15] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_17[15] <= Psram_Addr_To_Sram_FIFO_17[16];
        Psram_Addr_To_Sram_FIFO_18[15] <= Psram_Addr_To_Sram_FIFO_18[16];
        Psram_Addr_To_Sram_FIFO_19[15] <= Psram_Addr_To_Sram_FIFO_19[16];
        Psram_Addr_To_Sram_FIFO_20[15] <= Psram_Addr_To_Sram_FIFO_20[16];
        Psram_Addr_To_Sram_FIFO_21[15] <= Psram_Addr_To_Sram_FIFO_21[16];
        Psram_Addr_To_Sram_FIFO_22[15] <= Psram_Addr_To_Sram_FIFO_22[16];
        Psram_Addr_To_Sram_FIFO_23[15] <= Psram_Addr_To_Sram_FIFO_23[16];
        Psram_Addr_To_Sram_FIFO_24[15] <= Psram_Addr_To_Sram_FIFO_24[16];
        Psram_Addr_To_Sram_FIFO_25[15] <= Psram_Addr_To_Sram_FIFO_25[16];
        Psram_Addr_To_Sram_FIFO_26[15] <= Psram_Addr_To_Sram_FIFO_26[16];
        Psram_Addr_To_Sram_FIFO_27[15] <= Psram_Addr_To_Sram_FIFO_27[16];
        Psram_Addr_To_Sram_FIFO_28[15] <= Psram_Addr_To_Sram_FIFO_28[16];
        Psram_Addr_To_Sram_FIFO_29[15] <= Psram_Addr_To_Sram_FIFO_29[16];
        Psram_Addr_To_Sram_FIFO_30[15] <= Psram_Addr_To_Sram_FIFO_30[16];
        Psram_Addr_To_Sram_FIFO_31[15] <= Psram_Addr_To_Sram_FIFO_31[16];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_17[16] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_18[16] <= Psram_Addr_To_Sram_FIFO_18[17];
        Psram_Addr_To_Sram_FIFO_19[16] <= Psram_Addr_To_Sram_FIFO_19[17];
        Psram_Addr_To_Sram_FIFO_20[16] <= Psram_Addr_To_Sram_FIFO_20[17];
        Psram_Addr_To_Sram_FIFO_21[16] <= Psram_Addr_To_Sram_FIFO_21[17];
        Psram_Addr_To_Sram_FIFO_22[16] <= Psram_Addr_To_Sram_FIFO_22[17];
        Psram_Addr_To_Sram_FIFO_23[16] <= Psram_Addr_To_Sram_FIFO_23[17];
        Psram_Addr_To_Sram_FIFO_24[16] <= Psram_Addr_To_Sram_FIFO_24[17];
        Psram_Addr_To_Sram_FIFO_25[16] <= Psram_Addr_To_Sram_FIFO_25[17];
        Psram_Addr_To_Sram_FIFO_26[16] <= Psram_Addr_To_Sram_FIFO_26[17];
        Psram_Addr_To_Sram_FIFO_27[16] <= Psram_Addr_To_Sram_FIFO_27[17];
        Psram_Addr_To_Sram_FIFO_28[16] <= Psram_Addr_To_Sram_FIFO_28[17];
        Psram_Addr_To_Sram_FIFO_29[16] <= Psram_Addr_To_Sram_FIFO_29[17];
        Psram_Addr_To_Sram_FIFO_30[16] <= Psram_Addr_To_Sram_FIFO_30[17];
        Psram_Addr_To_Sram_FIFO_31[16] <= Psram_Addr_To_Sram_FIFO_31[17];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_18[17] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_19[17] <= Psram_Addr_To_Sram_FIFO_19[18];
        Psram_Addr_To_Sram_FIFO_20[17] <= Psram_Addr_To_Sram_FIFO_20[18];
        Psram_Addr_To_Sram_FIFO_21[17] <= Psram_Addr_To_Sram_FIFO_21[18];
        Psram_Addr_To_Sram_FIFO_22[17] <= Psram_Addr_To_Sram_FIFO_22[18];
        Psram_Addr_To_Sram_FIFO_23[17] <= Psram_Addr_To_Sram_FIFO_23[18];
        Psram_Addr_To_Sram_FIFO_24[17] <= Psram_Addr_To_Sram_FIFO_24[18];
        Psram_Addr_To_Sram_FIFO_25[17] <= Psram_Addr_To_Sram_FIFO_25[18];
        Psram_Addr_To_Sram_FIFO_26[17] <= Psram_Addr_To_Sram_FIFO_26[18];
        Psram_Addr_To_Sram_FIFO_27[17] <= Psram_Addr_To_Sram_FIFO_27[18];
        Psram_Addr_To_Sram_FIFO_28[17] <= Psram_Addr_To_Sram_FIFO_28[18];
        Psram_Addr_To_Sram_FIFO_29[17] <= Psram_Addr_To_Sram_FIFO_29[18];
        Psram_Addr_To_Sram_FIFO_30[17] <= Psram_Addr_To_Sram_FIFO_30[18];
        Psram_Addr_To_Sram_FIFO_31[17] <= Psram_Addr_To_Sram_FIFO_31[18];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_19[18] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_20[18] <= Psram_Addr_To_Sram_FIFO_20[19];
        Psram_Addr_To_Sram_FIFO_21[18] <= Psram_Addr_To_Sram_FIFO_21[19];
        Psram_Addr_To_Sram_FIFO_22[18] <= Psram_Addr_To_Sram_FIFO_22[19];
        Psram_Addr_To_Sram_FIFO_23[18] <= Psram_Addr_To_Sram_FIFO_23[19];
        Psram_Addr_To_Sram_FIFO_24[18] <= Psram_Addr_To_Sram_FIFO_24[19];
        Psram_Addr_To_Sram_FIFO_25[18] <= Psram_Addr_To_Sram_FIFO_25[19];
        Psram_Addr_To_Sram_FIFO_26[18] <= Psram_Addr_To_Sram_FIFO_26[19];
        Psram_Addr_To_Sram_FIFO_27[18] <= Psram_Addr_To_Sram_FIFO_27[19];
        Psram_Addr_To_Sram_FIFO_28[18] <= Psram_Addr_To_Sram_FIFO_28[19];
        Psram_Addr_To_Sram_FIFO_29[18] <= Psram_Addr_To_Sram_FIFO_29[19];
        Psram_Addr_To_Sram_FIFO_30[18] <= Psram_Addr_To_Sram_FIFO_30[19];
        Psram_Addr_To_Sram_FIFO_31[18] <= Psram_Addr_To_Sram_FIFO_31[19];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_20[19] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_21[19] <= Psram_Addr_To_Sram_FIFO_21[20];
        Psram_Addr_To_Sram_FIFO_22[19] <= Psram_Addr_To_Sram_FIFO_22[20];
        Psram_Addr_To_Sram_FIFO_23[19] <= Psram_Addr_To_Sram_FIFO_23[20];
        Psram_Addr_To_Sram_FIFO_24[19] <= Psram_Addr_To_Sram_FIFO_24[20];
        Psram_Addr_To_Sram_FIFO_25[19] <= Psram_Addr_To_Sram_FIFO_25[20];
        Psram_Addr_To_Sram_FIFO_26[19] <= Psram_Addr_To_Sram_FIFO_26[20];
        Psram_Addr_To_Sram_FIFO_27[19] <= Psram_Addr_To_Sram_FIFO_27[20];
        Psram_Addr_To_Sram_FIFO_28[19] <= Psram_Addr_To_Sram_FIFO_28[20];
        Psram_Addr_To_Sram_FIFO_29[19] <= Psram_Addr_To_Sram_FIFO_29[20];
        Psram_Addr_To_Sram_FIFO_30[19] <= Psram_Addr_To_Sram_FIFO_30[20];
        Psram_Addr_To_Sram_FIFO_31[19] <= Psram_Addr_To_Sram_FIFO_31[20];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_21[20] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_22[20] <= Psram_Addr_To_Sram_FIFO_22[21];
        Psram_Addr_To_Sram_FIFO_23[20] <= Psram_Addr_To_Sram_FIFO_23[21];
        Psram_Addr_To_Sram_FIFO_24[20] <= Psram_Addr_To_Sram_FIFO_24[21];
        Psram_Addr_To_Sram_FIFO_25[20] <= Psram_Addr_To_Sram_FIFO_25[21];
        Psram_Addr_To_Sram_FIFO_26[20] <= Psram_Addr_To_Sram_FIFO_26[21];
        Psram_Addr_To_Sram_FIFO_27[20] <= Psram_Addr_To_Sram_FIFO_27[21];
        Psram_Addr_To_Sram_FIFO_28[20] <= Psram_Addr_To_Sram_FIFO_28[21];
        Psram_Addr_To_Sram_FIFO_29[20] <= Psram_Addr_To_Sram_FIFO_29[21];
        Psram_Addr_To_Sram_FIFO_30[20] <= Psram_Addr_To_Sram_FIFO_30[21];
        Psram_Addr_To_Sram_FIFO_31[20] <= Psram_Addr_To_Sram_FIFO_31[21];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_22[21] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_23[21] <= Psram_Addr_To_Sram_FIFO_23[22];
        Psram_Addr_To_Sram_FIFO_24[21] <= Psram_Addr_To_Sram_FIFO_24[22];
        Psram_Addr_To_Sram_FIFO_25[21] <= Psram_Addr_To_Sram_FIFO_25[22];
        Psram_Addr_To_Sram_FIFO_26[21] <= Psram_Addr_To_Sram_FIFO_26[22];
        Psram_Addr_To_Sram_FIFO_27[21] <= Psram_Addr_To_Sram_FIFO_27[22];
        Psram_Addr_To_Sram_FIFO_28[21] <= Psram_Addr_To_Sram_FIFO_28[22];
        Psram_Addr_To_Sram_FIFO_29[21] <= Psram_Addr_To_Sram_FIFO_29[22];
        Psram_Addr_To_Sram_FIFO_30[21] <= Psram_Addr_To_Sram_FIFO_30[22];
        Psram_Addr_To_Sram_FIFO_31[21] <= Psram_Addr_To_Sram_FIFO_31[22];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_23[22] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_24[22] <= Psram_Addr_To_Sram_FIFO_24[23];
        Psram_Addr_To_Sram_FIFO_25[22] <= Psram_Addr_To_Sram_FIFO_25[23];
        Psram_Addr_To_Sram_FIFO_26[22] <= Psram_Addr_To_Sram_FIFO_26[23];
        Psram_Addr_To_Sram_FIFO_27[22] <= Psram_Addr_To_Sram_FIFO_27[23];
        Psram_Addr_To_Sram_FIFO_28[22] <= Psram_Addr_To_Sram_FIFO_28[23];
        Psram_Addr_To_Sram_FIFO_29[22] <= Psram_Addr_To_Sram_FIFO_29[23];
        Psram_Addr_To_Sram_FIFO_30[22] <= Psram_Addr_To_Sram_FIFO_30[23];
        Psram_Addr_To_Sram_FIFO_31[22] <= Psram_Addr_To_Sram_FIFO_31[23];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_24[23] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_25[23] <= Psram_Addr_To_Sram_FIFO_25[24];
        Psram_Addr_To_Sram_FIFO_26[23] <= Psram_Addr_To_Sram_FIFO_26[24];
        Psram_Addr_To_Sram_FIFO_27[23] <= Psram_Addr_To_Sram_FIFO_27[24];
        Psram_Addr_To_Sram_FIFO_28[23] <= Psram_Addr_To_Sram_FIFO_28[24];
        Psram_Addr_To_Sram_FIFO_29[23] <= Psram_Addr_To_Sram_FIFO_29[24];
        Psram_Addr_To_Sram_FIFO_30[23] <= Psram_Addr_To_Sram_FIFO_30[24];
        Psram_Addr_To_Sram_FIFO_31[23] <= Psram_Addr_To_Sram_FIFO_31[24];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_25[24] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_26[24] <= Psram_Addr_To_Sram_FIFO_26[25];
        Psram_Addr_To_Sram_FIFO_27[24] <= Psram_Addr_To_Sram_FIFO_27[25];
        Psram_Addr_To_Sram_FIFO_28[24] <= Psram_Addr_To_Sram_FIFO_28[25];
        Psram_Addr_To_Sram_FIFO_29[24] <= Psram_Addr_To_Sram_FIFO_29[25];
        Psram_Addr_To_Sram_FIFO_30[24] <= Psram_Addr_To_Sram_FIFO_30[25];
        Psram_Addr_To_Sram_FIFO_31[24] <= Psram_Addr_To_Sram_FIFO_31[25];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_26[25] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_27[25] <= Psram_Addr_To_Sram_FIFO_27[26];
        Psram_Addr_To_Sram_FIFO_28[25] <= Psram_Addr_To_Sram_FIFO_28[26];
        Psram_Addr_To_Sram_FIFO_29[25] <= Psram_Addr_To_Sram_FIFO_29[26];
        Psram_Addr_To_Sram_FIFO_30[25] <= Psram_Addr_To_Sram_FIFO_30[26];
        Psram_Addr_To_Sram_FIFO_31[25] <= Psram_Addr_To_Sram_FIFO_31[26];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_27[26] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_28[26] <= Psram_Addr_To_Sram_FIFO_28[27];
        Psram_Addr_To_Sram_FIFO_29[26] <= Psram_Addr_To_Sram_FIFO_29[27];
        Psram_Addr_To_Sram_FIFO_30[26] <= Psram_Addr_To_Sram_FIFO_30[27];
        Psram_Addr_To_Sram_FIFO_31[26] <= Psram_Addr_To_Sram_FIFO_31[27];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_28[27] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_29[27] <= Psram_Addr_To_Sram_FIFO_29[28];
        Psram_Addr_To_Sram_FIFO_30[27] <= Psram_Addr_To_Sram_FIFO_30[28];
        Psram_Addr_To_Sram_FIFO_31[27] <= Psram_Addr_To_Sram_FIFO_31[28];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_29[28] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_30[28] <= Psram_Addr_To_Sram_FIFO_30[29];
        Psram_Addr_To_Sram_FIFO_31[28] <= Psram_Addr_To_Sram_FIFO_31[29];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_30[29] <= i_Psram_Addr;
        Psram_Addr_To_Sram_FIFO_31[29] <= Psram_Addr_To_Sram_FIFO_31[30];
    end

    always @(posedge CLK) begin
        Psram_Addr_To_Sram_FIFO_31[30] <= i_Psram_Addr;
    end

    // Psram_En_To_Sram Logic
    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_1[0] <= i_Psram_En[1];
        Psram_En_To_Sram_FIFO_2[0] <= Psram_En_To_Sram_FIFO_2[1];
        Psram_En_To_Sram_FIFO_3[0] <= Psram_En_To_Sram_FIFO_3[1];
        Psram_En_To_Sram_FIFO_4[0] <= Psram_En_To_Sram_FIFO_4[1];
        Psram_En_To_Sram_FIFO_5[0] <= Psram_En_To_Sram_FIFO_5[1];
        Psram_En_To_Sram_FIFO_6[0] <= Psram_En_To_Sram_FIFO_6[1];
        Psram_En_To_Sram_FIFO_7[0] <= Psram_En_To_Sram_FIFO_7[1];
        Psram_En_To_Sram_FIFO_8[0] <= Psram_En_To_Sram_FIFO_8[1];
        Psram_En_To_Sram_FIFO_9[0] <= Psram_En_To_Sram_FIFO_9[1];
        Psram_En_To_Sram_FIFO_10[0] <= Psram_En_To_Sram_FIFO_10[1];
        Psram_En_To_Sram_FIFO_11[0] <= Psram_En_To_Sram_FIFO_11[1];
        Psram_En_To_Sram_FIFO_12[0] <= Psram_En_To_Sram_FIFO_12[1];
        Psram_En_To_Sram_FIFO_13[0] <= Psram_En_To_Sram_FIFO_13[1];
        Psram_En_To_Sram_FIFO_14[0] <= Psram_En_To_Sram_FIFO_14[1];
        Psram_En_To_Sram_FIFO_15[0] <= Psram_En_To_Sram_FIFO_15[1];
        Psram_En_To_Sram_FIFO_16[0] <= Psram_En_To_Sram_FIFO_16[1];
        Psram_En_To_Sram_FIFO_17[0] <= Psram_En_To_Sram_FIFO_17[1];
        Psram_En_To_Sram_FIFO_18[0] <= Psram_En_To_Sram_FIFO_18[1];
        Psram_En_To_Sram_FIFO_19[0] <= Psram_En_To_Sram_FIFO_19[1];
        Psram_En_To_Sram_FIFO_20[0] <= Psram_En_To_Sram_FIFO_20[1];
        Psram_En_To_Sram_FIFO_21[0] <= Psram_En_To_Sram_FIFO_21[1];
        Psram_En_To_Sram_FIFO_22[0] <= Psram_En_To_Sram_FIFO_22[1];
        Psram_En_To_Sram_FIFO_23[0] <= Psram_En_To_Sram_FIFO_23[1];
        Psram_En_To_Sram_FIFO_24[0] <= Psram_En_To_Sram_FIFO_24[1];
        Psram_En_To_Sram_FIFO_25[0] <= Psram_En_To_Sram_FIFO_25[1];
        Psram_En_To_Sram_FIFO_26[0] <= Psram_En_To_Sram_FIFO_26[1];
        Psram_En_To_Sram_FIFO_27[0] <= Psram_En_To_Sram_FIFO_27[1];
        Psram_En_To_Sram_FIFO_28[0] <= Psram_En_To_Sram_FIFO_28[1];
        Psram_En_To_Sram_FIFO_29[0] <= Psram_En_To_Sram_FIFO_29[1];
        Psram_En_To_Sram_FIFO_30[0] <= Psram_En_To_Sram_FIFO_30[1];
        Psram_En_To_Sram_FIFO_31[0] <= Psram_En_To_Sram_FIFO_31[1];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_2[1] <= i_Psram_En[2];
        Psram_En_To_Sram_FIFO_3[1] <= Psram_En_To_Sram_FIFO_3[2];
        Psram_En_To_Sram_FIFO_4[1] <= Psram_En_To_Sram_FIFO_4[2];
        Psram_En_To_Sram_FIFO_5[1] <= Psram_En_To_Sram_FIFO_5[2];
        Psram_En_To_Sram_FIFO_6[1] <= Psram_En_To_Sram_FIFO_6[2];
        Psram_En_To_Sram_FIFO_7[1] <= Psram_En_To_Sram_FIFO_7[2];
        Psram_En_To_Sram_FIFO_8[1] <= Psram_En_To_Sram_FIFO_8[2];
        Psram_En_To_Sram_FIFO_9[1] <= Psram_En_To_Sram_FIFO_9[2];
        Psram_En_To_Sram_FIFO_10[1] <= Psram_En_To_Sram_FIFO_10[2];
        Psram_En_To_Sram_FIFO_11[1] <= Psram_En_To_Sram_FIFO_11[2];
        Psram_En_To_Sram_FIFO_12[1] <= Psram_En_To_Sram_FIFO_12[2];
        Psram_En_To_Sram_FIFO_13[1] <= Psram_En_To_Sram_FIFO_13[2];
        Psram_En_To_Sram_FIFO_14[1] <= Psram_En_To_Sram_FIFO_14[2];
        Psram_En_To_Sram_FIFO_15[1] <= Psram_En_To_Sram_FIFO_15[2];
        Psram_En_To_Sram_FIFO_16[1] <= Psram_En_To_Sram_FIFO_16[2];
        Psram_En_To_Sram_FIFO_17[1] <= Psram_En_To_Sram_FIFO_17[2];
        Psram_En_To_Sram_FIFO_18[1] <= Psram_En_To_Sram_FIFO_18[2];
        Psram_En_To_Sram_FIFO_19[1] <= Psram_En_To_Sram_FIFO_19[2];
        Psram_En_To_Sram_FIFO_20[1] <= Psram_En_To_Sram_FIFO_20[2];
        Psram_En_To_Sram_FIFO_21[1] <= Psram_En_To_Sram_FIFO_21[2];
        Psram_En_To_Sram_FIFO_22[1] <= Psram_En_To_Sram_FIFO_22[2];
        Psram_En_To_Sram_FIFO_23[1] <= Psram_En_To_Sram_FIFO_23[2];
        Psram_En_To_Sram_FIFO_24[1] <= Psram_En_To_Sram_FIFO_24[2];
        Psram_En_To_Sram_FIFO_25[1] <= Psram_En_To_Sram_FIFO_25[2];
        Psram_En_To_Sram_FIFO_26[1] <= Psram_En_To_Sram_FIFO_26[2];
        Psram_En_To_Sram_FIFO_27[1] <= Psram_En_To_Sram_FIFO_27[2];
        Psram_En_To_Sram_FIFO_28[1] <= Psram_En_To_Sram_FIFO_28[2];
        Psram_En_To_Sram_FIFO_29[1] <= Psram_En_To_Sram_FIFO_29[2];
        Psram_En_To_Sram_FIFO_30[1] <= Psram_En_To_Sram_FIFO_30[2];
        Psram_En_To_Sram_FIFO_31[1] <= Psram_En_To_Sram_FIFO_31[2];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_3[2] <= i_Psram_En[3];
        Psram_En_To_Sram_FIFO_4[2] <= Psram_En_To_Sram_FIFO_4[3];
        Psram_En_To_Sram_FIFO_5[2] <= Psram_En_To_Sram_FIFO_5[3];
        Psram_En_To_Sram_FIFO_6[2] <= Psram_En_To_Sram_FIFO_6[3];
        Psram_En_To_Sram_FIFO_7[2] <= Psram_En_To_Sram_FIFO_7[3];
        Psram_En_To_Sram_FIFO_8[2] <= Psram_En_To_Sram_FIFO_8[3];
        Psram_En_To_Sram_FIFO_9[2] <= Psram_En_To_Sram_FIFO_9[3];
        Psram_En_To_Sram_FIFO_10[2] <= Psram_En_To_Sram_FIFO_10[3];
        Psram_En_To_Sram_FIFO_11[2] <= Psram_En_To_Sram_FIFO_11[3];
        Psram_En_To_Sram_FIFO_12[2] <= Psram_En_To_Sram_FIFO_12[3];
        Psram_En_To_Sram_FIFO_13[2] <= Psram_En_To_Sram_FIFO_13[3];
        Psram_En_To_Sram_FIFO_14[2] <= Psram_En_To_Sram_FIFO_14[3];
        Psram_En_To_Sram_FIFO_15[2] <= Psram_En_To_Sram_FIFO_15[3];
        Psram_En_To_Sram_FIFO_16[2] <= Psram_En_To_Sram_FIFO_16[3];
        Psram_En_To_Sram_FIFO_17[2] <= Psram_En_To_Sram_FIFO_17[3];
        Psram_En_To_Sram_FIFO_18[2] <= Psram_En_To_Sram_FIFO_18[3];
        Psram_En_To_Sram_FIFO_19[2] <= Psram_En_To_Sram_FIFO_19[3];
        Psram_En_To_Sram_FIFO_20[2] <= Psram_En_To_Sram_FIFO_20[3];
        Psram_En_To_Sram_FIFO_21[2] <= Psram_En_To_Sram_FIFO_21[3];
        Psram_En_To_Sram_FIFO_22[2] <= Psram_En_To_Sram_FIFO_22[3];
        Psram_En_To_Sram_FIFO_23[2] <= Psram_En_To_Sram_FIFO_23[3];
        Psram_En_To_Sram_FIFO_24[2] <= Psram_En_To_Sram_FIFO_24[3];
        Psram_En_To_Sram_FIFO_25[2] <= Psram_En_To_Sram_FIFO_25[3];
        Psram_En_To_Sram_FIFO_26[2] <= Psram_En_To_Sram_FIFO_26[3];
        Psram_En_To_Sram_FIFO_27[2] <= Psram_En_To_Sram_FIFO_27[3];
        Psram_En_To_Sram_FIFO_28[2] <= Psram_En_To_Sram_FIFO_28[3];
        Psram_En_To_Sram_FIFO_29[2] <= Psram_En_To_Sram_FIFO_29[3];
        Psram_En_To_Sram_FIFO_30[2] <= Psram_En_To_Sram_FIFO_30[3];
        Psram_En_To_Sram_FIFO_31[2] <= Psram_En_To_Sram_FIFO_31[3];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_4[3] <= i_Psram_En[4];
        Psram_En_To_Sram_FIFO_5[3] <= Psram_En_To_Sram_FIFO_5[4];
        Psram_En_To_Sram_FIFO_6[3] <= Psram_En_To_Sram_FIFO_6[4];
        Psram_En_To_Sram_FIFO_7[3] <= Psram_En_To_Sram_FIFO_7[4];
        Psram_En_To_Sram_FIFO_8[3] <= Psram_En_To_Sram_FIFO_8[4];
        Psram_En_To_Sram_FIFO_9[3] <= Psram_En_To_Sram_FIFO_9[4];
        Psram_En_To_Sram_FIFO_10[3] <= Psram_En_To_Sram_FIFO_10[4];
        Psram_En_To_Sram_FIFO_11[3] <= Psram_En_To_Sram_FIFO_11[4];
        Psram_En_To_Sram_FIFO_12[3] <= Psram_En_To_Sram_FIFO_12[4];
        Psram_En_To_Sram_FIFO_13[3] <= Psram_En_To_Sram_FIFO_13[4];
        Psram_En_To_Sram_FIFO_14[3] <= Psram_En_To_Sram_FIFO_14[4];
        Psram_En_To_Sram_FIFO_15[3] <= Psram_En_To_Sram_FIFO_15[4];
        Psram_En_To_Sram_FIFO_16[3] <= Psram_En_To_Sram_FIFO_16[4];
        Psram_En_To_Sram_FIFO_17[3] <= Psram_En_To_Sram_FIFO_17[4];
        Psram_En_To_Sram_FIFO_18[3] <= Psram_En_To_Sram_FIFO_18[4];
        Psram_En_To_Sram_FIFO_19[3] <= Psram_En_To_Sram_FIFO_19[4];
        Psram_En_To_Sram_FIFO_20[3] <= Psram_En_To_Sram_FIFO_20[4];
        Psram_En_To_Sram_FIFO_21[3] <= Psram_En_To_Sram_FIFO_21[4];
        Psram_En_To_Sram_FIFO_22[3] <= Psram_En_To_Sram_FIFO_22[4];
        Psram_En_To_Sram_FIFO_23[3] <= Psram_En_To_Sram_FIFO_23[4];
        Psram_En_To_Sram_FIFO_24[3] <= Psram_En_To_Sram_FIFO_24[4];
        Psram_En_To_Sram_FIFO_25[3] <= Psram_En_To_Sram_FIFO_25[4];
        Psram_En_To_Sram_FIFO_26[3] <= Psram_En_To_Sram_FIFO_26[4];
        Psram_En_To_Sram_FIFO_27[3] <= Psram_En_To_Sram_FIFO_27[4];
        Psram_En_To_Sram_FIFO_28[3] <= Psram_En_To_Sram_FIFO_28[4];
        Psram_En_To_Sram_FIFO_29[3] <= Psram_En_To_Sram_FIFO_29[4];
        Psram_En_To_Sram_FIFO_30[3] <= Psram_En_To_Sram_FIFO_30[4];
        Psram_En_To_Sram_FIFO_31[3] <= Psram_En_To_Sram_FIFO_31[4];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_5[4] <= i_Psram_En[5];
        Psram_En_To_Sram_FIFO_6[4] <= Psram_En_To_Sram_FIFO_6[5];
        Psram_En_To_Sram_FIFO_7[4] <= Psram_En_To_Sram_FIFO_7[5];
        Psram_En_To_Sram_FIFO_8[4] <= Psram_En_To_Sram_FIFO_8[5];
        Psram_En_To_Sram_FIFO_9[4] <= Psram_En_To_Sram_FIFO_9[5];
        Psram_En_To_Sram_FIFO_10[4] <= Psram_En_To_Sram_FIFO_10[5];
        Psram_En_To_Sram_FIFO_11[4] <= Psram_En_To_Sram_FIFO_11[5];
        Psram_En_To_Sram_FIFO_12[4] <= Psram_En_To_Sram_FIFO_12[5];
        Psram_En_To_Sram_FIFO_13[4] <= Psram_En_To_Sram_FIFO_13[5];
        Psram_En_To_Sram_FIFO_14[4] <= Psram_En_To_Sram_FIFO_14[5];
        Psram_En_To_Sram_FIFO_15[4] <= Psram_En_To_Sram_FIFO_15[5];
        Psram_En_To_Sram_FIFO_16[4] <= Psram_En_To_Sram_FIFO_16[5];
        Psram_En_To_Sram_FIFO_17[4] <= Psram_En_To_Sram_FIFO_17[5];
        Psram_En_To_Sram_FIFO_18[4] <= Psram_En_To_Sram_FIFO_18[5];
        Psram_En_To_Sram_FIFO_19[4] <= Psram_En_To_Sram_FIFO_19[5];
        Psram_En_To_Sram_FIFO_20[4] <= Psram_En_To_Sram_FIFO_20[5];
        Psram_En_To_Sram_FIFO_21[4] <= Psram_En_To_Sram_FIFO_21[5];
        Psram_En_To_Sram_FIFO_22[4] <= Psram_En_To_Sram_FIFO_22[5];
        Psram_En_To_Sram_FIFO_23[4] <= Psram_En_To_Sram_FIFO_23[5];
        Psram_En_To_Sram_FIFO_24[4] <= Psram_En_To_Sram_FIFO_24[5];
        Psram_En_To_Sram_FIFO_25[4] <= Psram_En_To_Sram_FIFO_25[5];
        Psram_En_To_Sram_FIFO_26[4] <= Psram_En_To_Sram_FIFO_26[5];
        Psram_En_To_Sram_FIFO_27[4] <= Psram_En_To_Sram_FIFO_27[5];
        Psram_En_To_Sram_FIFO_28[4] <= Psram_En_To_Sram_FIFO_28[5];
        Psram_En_To_Sram_FIFO_29[4] <= Psram_En_To_Sram_FIFO_29[5];
        Psram_En_To_Sram_FIFO_30[4] <= Psram_En_To_Sram_FIFO_30[5];
        Psram_En_To_Sram_FIFO_31[4] <= Psram_En_To_Sram_FIFO_31[5];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_6[5] <= i_Psram_En[6];
        Psram_En_To_Sram_FIFO_7[5] <= Psram_En_To_Sram_FIFO_7[6];
        Psram_En_To_Sram_FIFO_8[5] <= Psram_En_To_Sram_FIFO_8[6];
        Psram_En_To_Sram_FIFO_9[5] <= Psram_En_To_Sram_FIFO_9[6];
        Psram_En_To_Sram_FIFO_10[5] <= Psram_En_To_Sram_FIFO_10[6];
        Psram_En_To_Sram_FIFO_11[5] <= Psram_En_To_Sram_FIFO_11[6];
        Psram_En_To_Sram_FIFO_12[5] <= Psram_En_To_Sram_FIFO_12[6];
        Psram_En_To_Sram_FIFO_13[5] <= Psram_En_To_Sram_FIFO_13[6];
        Psram_En_To_Sram_FIFO_14[5] <= Psram_En_To_Sram_FIFO_14[6];
        Psram_En_To_Sram_FIFO_15[5] <= Psram_En_To_Sram_FIFO_15[6];
        Psram_En_To_Sram_FIFO_16[5] <= Psram_En_To_Sram_FIFO_16[6];
        Psram_En_To_Sram_FIFO_17[5] <= Psram_En_To_Sram_FIFO_17[6];
        Psram_En_To_Sram_FIFO_18[5] <= Psram_En_To_Sram_FIFO_18[6];
        Psram_En_To_Sram_FIFO_19[5] <= Psram_En_To_Sram_FIFO_19[6];
        Psram_En_To_Sram_FIFO_20[5] <= Psram_En_To_Sram_FIFO_20[6];
        Psram_En_To_Sram_FIFO_21[5] <= Psram_En_To_Sram_FIFO_21[6];
        Psram_En_To_Sram_FIFO_22[5] <= Psram_En_To_Sram_FIFO_22[6];
        Psram_En_To_Sram_FIFO_23[5] <= Psram_En_To_Sram_FIFO_23[6];
        Psram_En_To_Sram_FIFO_24[5] <= Psram_En_To_Sram_FIFO_24[6];
        Psram_En_To_Sram_FIFO_25[5] <= Psram_En_To_Sram_FIFO_25[6];
        Psram_En_To_Sram_FIFO_26[5] <= Psram_En_To_Sram_FIFO_26[6];
        Psram_En_To_Sram_FIFO_27[5] <= Psram_En_To_Sram_FIFO_27[6];
        Psram_En_To_Sram_FIFO_28[5] <= Psram_En_To_Sram_FIFO_28[6];
        Psram_En_To_Sram_FIFO_29[5] <= Psram_En_To_Sram_FIFO_29[6];
        Psram_En_To_Sram_FIFO_30[5] <= Psram_En_To_Sram_FIFO_30[6];
        Psram_En_To_Sram_FIFO_31[5] <= Psram_En_To_Sram_FIFO_31[6];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_7[6] <= i_Psram_En[7];
        Psram_En_To_Sram_FIFO_8[6] <= Psram_En_To_Sram_FIFO_8[7];
        Psram_En_To_Sram_FIFO_9[6] <= Psram_En_To_Sram_FIFO_9[7];
        Psram_En_To_Sram_FIFO_10[6] <= Psram_En_To_Sram_FIFO_10[7];
        Psram_En_To_Sram_FIFO_11[6] <= Psram_En_To_Sram_FIFO_11[7];
        Psram_En_To_Sram_FIFO_12[6] <= Psram_En_To_Sram_FIFO_12[7];
        Psram_En_To_Sram_FIFO_13[6] <= Psram_En_To_Sram_FIFO_13[7];
        Psram_En_To_Sram_FIFO_14[6] <= Psram_En_To_Sram_FIFO_14[7];
        Psram_En_To_Sram_FIFO_15[6] <= Psram_En_To_Sram_FIFO_15[7];
        Psram_En_To_Sram_FIFO_16[6] <= Psram_En_To_Sram_FIFO_16[7];
        Psram_En_To_Sram_FIFO_17[6] <= Psram_En_To_Sram_FIFO_17[7];
        Psram_En_To_Sram_FIFO_18[6] <= Psram_En_To_Sram_FIFO_18[7];
        Psram_En_To_Sram_FIFO_19[6] <= Psram_En_To_Sram_FIFO_19[7];
        Psram_En_To_Sram_FIFO_20[6] <= Psram_En_To_Sram_FIFO_20[7];
        Psram_En_To_Sram_FIFO_21[6] <= Psram_En_To_Sram_FIFO_21[7];
        Psram_En_To_Sram_FIFO_22[6] <= Psram_En_To_Sram_FIFO_22[7];
        Psram_En_To_Sram_FIFO_23[6] <= Psram_En_To_Sram_FIFO_23[7];
        Psram_En_To_Sram_FIFO_24[6] <= Psram_En_To_Sram_FIFO_24[7];
        Psram_En_To_Sram_FIFO_25[6] <= Psram_En_To_Sram_FIFO_25[7];
        Psram_En_To_Sram_FIFO_26[6] <= Psram_En_To_Sram_FIFO_26[7];
        Psram_En_To_Sram_FIFO_27[6] <= Psram_En_To_Sram_FIFO_27[7];
        Psram_En_To_Sram_FIFO_28[6] <= Psram_En_To_Sram_FIFO_28[7];
        Psram_En_To_Sram_FIFO_29[6] <= Psram_En_To_Sram_FIFO_29[7];
        Psram_En_To_Sram_FIFO_30[6] <= Psram_En_To_Sram_FIFO_30[7];
        Psram_En_To_Sram_FIFO_31[6] <= Psram_En_To_Sram_FIFO_31[7];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_8[7] <= i_Psram_En[8];
        Psram_En_To_Sram_FIFO_9[7] <= Psram_En_To_Sram_FIFO_9[8];
        Psram_En_To_Sram_FIFO_10[7] <= Psram_En_To_Sram_FIFO_10[8];
        Psram_En_To_Sram_FIFO_11[7] <= Psram_En_To_Sram_FIFO_11[8];
        Psram_En_To_Sram_FIFO_12[7] <= Psram_En_To_Sram_FIFO_12[8];
        Psram_En_To_Sram_FIFO_13[7] <= Psram_En_To_Sram_FIFO_13[8];
        Psram_En_To_Sram_FIFO_14[7] <= Psram_En_To_Sram_FIFO_14[8];
        Psram_En_To_Sram_FIFO_15[7] <= Psram_En_To_Sram_FIFO_15[8];
        Psram_En_To_Sram_FIFO_16[7] <= Psram_En_To_Sram_FIFO_16[8];
        Psram_En_To_Sram_FIFO_17[7] <= Psram_En_To_Sram_FIFO_17[8];
        Psram_En_To_Sram_FIFO_18[7] <= Psram_En_To_Sram_FIFO_18[8];
        Psram_En_To_Sram_FIFO_19[7] <= Psram_En_To_Sram_FIFO_19[8];
        Psram_En_To_Sram_FIFO_20[7] <= Psram_En_To_Sram_FIFO_20[8];
        Psram_En_To_Sram_FIFO_21[7] <= Psram_En_To_Sram_FIFO_21[8];
        Psram_En_To_Sram_FIFO_22[7] <= Psram_En_To_Sram_FIFO_22[8];
        Psram_En_To_Sram_FIFO_23[7] <= Psram_En_To_Sram_FIFO_23[8];
        Psram_En_To_Sram_FIFO_24[7] <= Psram_En_To_Sram_FIFO_24[8];
        Psram_En_To_Sram_FIFO_25[7] <= Psram_En_To_Sram_FIFO_25[8];
        Psram_En_To_Sram_FIFO_26[7] <= Psram_En_To_Sram_FIFO_26[8];
        Psram_En_To_Sram_FIFO_27[7] <= Psram_En_To_Sram_FIFO_27[8];
        Psram_En_To_Sram_FIFO_28[7] <= Psram_En_To_Sram_FIFO_28[8];
        Psram_En_To_Sram_FIFO_29[7] <= Psram_En_To_Sram_FIFO_29[8];
        Psram_En_To_Sram_FIFO_30[7] <= Psram_En_To_Sram_FIFO_30[8];
        Psram_En_To_Sram_FIFO_31[7] <= Psram_En_To_Sram_FIFO_31[8];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_9[8] <= i_Psram_En[9];
        Psram_En_To_Sram_FIFO_10[8] <= Psram_En_To_Sram_FIFO_10[9];
        Psram_En_To_Sram_FIFO_11[8] <= Psram_En_To_Sram_FIFO_11[9];
        Psram_En_To_Sram_FIFO_12[8] <= Psram_En_To_Sram_FIFO_12[9];
        Psram_En_To_Sram_FIFO_13[8] <= Psram_En_To_Sram_FIFO_13[9];
        Psram_En_To_Sram_FIFO_14[8] <= Psram_En_To_Sram_FIFO_14[9];
        Psram_En_To_Sram_FIFO_15[8] <= Psram_En_To_Sram_FIFO_15[9];
        Psram_En_To_Sram_FIFO_16[8] <= Psram_En_To_Sram_FIFO_16[9];
        Psram_En_To_Sram_FIFO_17[8] <= Psram_En_To_Sram_FIFO_17[9];
        Psram_En_To_Sram_FIFO_18[8] <= Psram_En_To_Sram_FIFO_18[9];
        Psram_En_To_Sram_FIFO_19[8] <= Psram_En_To_Sram_FIFO_19[9];
        Psram_En_To_Sram_FIFO_20[8] <= Psram_En_To_Sram_FIFO_20[9];
        Psram_En_To_Sram_FIFO_21[8] <= Psram_En_To_Sram_FIFO_21[9];
        Psram_En_To_Sram_FIFO_22[8] <= Psram_En_To_Sram_FIFO_22[9];
        Psram_En_To_Sram_FIFO_23[8] <= Psram_En_To_Sram_FIFO_23[9];
        Psram_En_To_Sram_FIFO_24[8] <= Psram_En_To_Sram_FIFO_24[9];
        Psram_En_To_Sram_FIFO_25[8] <= Psram_En_To_Sram_FIFO_25[9];
        Psram_En_To_Sram_FIFO_26[8] <= Psram_En_To_Sram_FIFO_26[9];
        Psram_En_To_Sram_FIFO_27[8] <= Psram_En_To_Sram_FIFO_27[9];
        Psram_En_To_Sram_FIFO_28[8] <= Psram_En_To_Sram_FIFO_28[9];
        Psram_En_To_Sram_FIFO_29[8] <= Psram_En_To_Sram_FIFO_29[9];
        Psram_En_To_Sram_FIFO_30[8] <= Psram_En_To_Sram_FIFO_30[9];
        Psram_En_To_Sram_FIFO_31[8] <= Psram_En_To_Sram_FIFO_31[9];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_10[9] <= i_Psram_En[10];
        Psram_En_To_Sram_FIFO_11[9] <= Psram_En_To_Sram_FIFO_11[10];
        Psram_En_To_Sram_FIFO_12[9] <= Psram_En_To_Sram_FIFO_12[10];
        Psram_En_To_Sram_FIFO_13[9] <= Psram_En_To_Sram_FIFO_13[10];
        Psram_En_To_Sram_FIFO_14[9] <= Psram_En_To_Sram_FIFO_14[10];
        Psram_En_To_Sram_FIFO_15[9] <= Psram_En_To_Sram_FIFO_15[10];
        Psram_En_To_Sram_FIFO_16[9] <= Psram_En_To_Sram_FIFO_16[10];
        Psram_En_To_Sram_FIFO_17[9] <= Psram_En_To_Sram_FIFO_17[10];
        Psram_En_To_Sram_FIFO_18[9] <= Psram_En_To_Sram_FIFO_18[10];
        Psram_En_To_Sram_FIFO_19[9] <= Psram_En_To_Sram_FIFO_19[10];
        Psram_En_To_Sram_FIFO_20[9] <= Psram_En_To_Sram_FIFO_20[10];
        Psram_En_To_Sram_FIFO_21[9] <= Psram_En_To_Sram_FIFO_21[10];
        Psram_En_To_Sram_FIFO_22[9] <= Psram_En_To_Sram_FIFO_22[10];
        Psram_En_To_Sram_FIFO_23[9] <= Psram_En_To_Sram_FIFO_23[10];
        Psram_En_To_Sram_FIFO_24[9] <= Psram_En_To_Sram_FIFO_24[10];
        Psram_En_To_Sram_FIFO_25[9] <= Psram_En_To_Sram_FIFO_25[10];
        Psram_En_To_Sram_FIFO_26[9] <= Psram_En_To_Sram_FIFO_26[10];
        Psram_En_To_Sram_FIFO_27[9] <= Psram_En_To_Sram_FIFO_27[10];
        Psram_En_To_Sram_FIFO_28[9] <= Psram_En_To_Sram_FIFO_28[10];
        Psram_En_To_Sram_FIFO_29[9] <= Psram_En_To_Sram_FIFO_29[10];
        Psram_En_To_Sram_FIFO_30[9] <= Psram_En_To_Sram_FIFO_30[10];
        Psram_En_To_Sram_FIFO_31[9] <= Psram_En_To_Sram_FIFO_31[10];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_11[10] <= i_Psram_En[11];
        Psram_En_To_Sram_FIFO_12[10] <= Psram_En_To_Sram_FIFO_12[11];
        Psram_En_To_Sram_FIFO_13[10] <= Psram_En_To_Sram_FIFO_13[11];
        Psram_En_To_Sram_FIFO_14[10] <= Psram_En_To_Sram_FIFO_14[11];
        Psram_En_To_Sram_FIFO_15[10] <= Psram_En_To_Sram_FIFO_15[11];
        Psram_En_To_Sram_FIFO_16[10] <= Psram_En_To_Sram_FIFO_16[11];
        Psram_En_To_Sram_FIFO_17[10] <= Psram_En_To_Sram_FIFO_17[11];
        Psram_En_To_Sram_FIFO_18[10] <= Psram_En_To_Sram_FIFO_18[11];
        Psram_En_To_Sram_FIFO_19[10] <= Psram_En_To_Sram_FIFO_19[11];
        Psram_En_To_Sram_FIFO_20[10] <= Psram_En_To_Sram_FIFO_20[11];
        Psram_En_To_Sram_FIFO_21[10] <= Psram_En_To_Sram_FIFO_21[11];
        Psram_En_To_Sram_FIFO_22[10] <= Psram_En_To_Sram_FIFO_22[11];
        Psram_En_To_Sram_FIFO_23[10] <= Psram_En_To_Sram_FIFO_23[11];
        Psram_En_To_Sram_FIFO_24[10] <= Psram_En_To_Sram_FIFO_24[11];
        Psram_En_To_Sram_FIFO_25[10] <= Psram_En_To_Sram_FIFO_25[11];
        Psram_En_To_Sram_FIFO_26[10] <= Psram_En_To_Sram_FIFO_26[11];
        Psram_En_To_Sram_FIFO_27[10] <= Psram_En_To_Sram_FIFO_27[11];
        Psram_En_To_Sram_FIFO_28[10] <= Psram_En_To_Sram_FIFO_28[11];
        Psram_En_To_Sram_FIFO_29[10] <= Psram_En_To_Sram_FIFO_29[11];
        Psram_En_To_Sram_FIFO_30[10] <= Psram_En_To_Sram_FIFO_30[11];
        Psram_En_To_Sram_FIFO_31[10] <= Psram_En_To_Sram_FIFO_31[11];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_12[11] <= i_Psram_En[12];
        Psram_En_To_Sram_FIFO_13[11] <= Psram_En_To_Sram_FIFO_13[12];
        Psram_En_To_Sram_FIFO_14[11] <= Psram_En_To_Sram_FIFO_14[12];
        Psram_En_To_Sram_FIFO_15[11] <= Psram_En_To_Sram_FIFO_15[12];
        Psram_En_To_Sram_FIFO_16[11] <= Psram_En_To_Sram_FIFO_16[12];
        Psram_En_To_Sram_FIFO_17[11] <= Psram_En_To_Sram_FIFO_17[12];
        Psram_En_To_Sram_FIFO_18[11] <= Psram_En_To_Sram_FIFO_18[12];
        Psram_En_To_Sram_FIFO_19[11] <= Psram_En_To_Sram_FIFO_19[12];
        Psram_En_To_Sram_FIFO_20[11] <= Psram_En_To_Sram_FIFO_20[12];
        Psram_En_To_Sram_FIFO_21[11] <= Psram_En_To_Sram_FIFO_21[12];
        Psram_En_To_Sram_FIFO_22[11] <= Psram_En_To_Sram_FIFO_22[12];
        Psram_En_To_Sram_FIFO_23[11] <= Psram_En_To_Sram_FIFO_23[12];
        Psram_En_To_Sram_FIFO_24[11] <= Psram_En_To_Sram_FIFO_24[12];
        Psram_En_To_Sram_FIFO_25[11] <= Psram_En_To_Sram_FIFO_25[12];
        Psram_En_To_Sram_FIFO_26[11] <= Psram_En_To_Sram_FIFO_26[12];
        Psram_En_To_Sram_FIFO_27[11] <= Psram_En_To_Sram_FIFO_27[12];
        Psram_En_To_Sram_FIFO_28[11] <= Psram_En_To_Sram_FIFO_28[12];
        Psram_En_To_Sram_FIFO_29[11] <= Psram_En_To_Sram_FIFO_29[12];
        Psram_En_To_Sram_FIFO_30[11] <= Psram_En_To_Sram_FIFO_30[12];
        Psram_En_To_Sram_FIFO_31[11] <= Psram_En_To_Sram_FIFO_31[12];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_13[12] <= i_Psram_En[13];
        Psram_En_To_Sram_FIFO_14[12] <= Psram_En_To_Sram_FIFO_14[13];
        Psram_En_To_Sram_FIFO_15[12] <= Psram_En_To_Sram_FIFO_15[13];
        Psram_En_To_Sram_FIFO_16[12] <= Psram_En_To_Sram_FIFO_16[13];
        Psram_En_To_Sram_FIFO_17[12] <= Psram_En_To_Sram_FIFO_17[13];
        Psram_En_To_Sram_FIFO_18[12] <= Psram_En_To_Sram_FIFO_18[13];
        Psram_En_To_Sram_FIFO_19[12] <= Psram_En_To_Sram_FIFO_19[13];
        Psram_En_To_Sram_FIFO_20[12] <= Psram_En_To_Sram_FIFO_20[13];
        Psram_En_To_Sram_FIFO_21[12] <= Psram_En_To_Sram_FIFO_21[13];
        Psram_En_To_Sram_FIFO_22[12] <= Psram_En_To_Sram_FIFO_22[13];
        Psram_En_To_Sram_FIFO_23[12] <= Psram_En_To_Sram_FIFO_23[13];
        Psram_En_To_Sram_FIFO_24[12] <= Psram_En_To_Sram_FIFO_24[13];
        Psram_En_To_Sram_FIFO_25[12] <= Psram_En_To_Sram_FIFO_25[13];
        Psram_En_To_Sram_FIFO_26[12] <= Psram_En_To_Sram_FIFO_26[13];
        Psram_En_To_Sram_FIFO_27[12] <= Psram_En_To_Sram_FIFO_27[13];
        Psram_En_To_Sram_FIFO_28[12] <= Psram_En_To_Sram_FIFO_28[13];
        Psram_En_To_Sram_FIFO_29[12] <= Psram_En_To_Sram_FIFO_29[13];
        Psram_En_To_Sram_FIFO_30[12] <= Psram_En_To_Sram_FIFO_30[13];
        Psram_En_To_Sram_FIFO_31[12] <= Psram_En_To_Sram_FIFO_31[13];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_14[13] <= i_Psram_En[14];
        Psram_En_To_Sram_FIFO_15[13] <= Psram_En_To_Sram_FIFO_15[14];
        Psram_En_To_Sram_FIFO_16[13] <= Psram_En_To_Sram_FIFO_16[14];
        Psram_En_To_Sram_FIFO_17[13] <= Psram_En_To_Sram_FIFO_17[14];
        Psram_En_To_Sram_FIFO_18[13] <= Psram_En_To_Sram_FIFO_18[14];
        Psram_En_To_Sram_FIFO_19[13] <= Psram_En_To_Sram_FIFO_19[14];
        Psram_En_To_Sram_FIFO_20[13] <= Psram_En_To_Sram_FIFO_20[14];
        Psram_En_To_Sram_FIFO_21[13] <= Psram_En_To_Sram_FIFO_21[14];
        Psram_En_To_Sram_FIFO_22[13] <= Psram_En_To_Sram_FIFO_22[14];
        Psram_En_To_Sram_FIFO_23[13] <= Psram_En_To_Sram_FIFO_23[14];
        Psram_En_To_Sram_FIFO_24[13] <= Psram_En_To_Sram_FIFO_24[14];
        Psram_En_To_Sram_FIFO_25[13] <= Psram_En_To_Sram_FIFO_25[14];
        Psram_En_To_Sram_FIFO_26[13] <= Psram_En_To_Sram_FIFO_26[14];
        Psram_En_To_Sram_FIFO_27[13] <= Psram_En_To_Sram_FIFO_27[14];
        Psram_En_To_Sram_FIFO_28[13] <= Psram_En_To_Sram_FIFO_28[14];
        Psram_En_To_Sram_FIFO_29[13] <= Psram_En_To_Sram_FIFO_29[14];
        Psram_En_To_Sram_FIFO_30[13] <= Psram_En_To_Sram_FIFO_30[14];
        Psram_En_To_Sram_FIFO_31[13] <= Psram_En_To_Sram_FIFO_31[14];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_15[14] <= i_Psram_En[15];
        Psram_En_To_Sram_FIFO_16[14] <= Psram_En_To_Sram_FIFO_16[15];
        Psram_En_To_Sram_FIFO_17[14] <= Psram_En_To_Sram_FIFO_17[15];
        Psram_En_To_Sram_FIFO_18[14] <= Psram_En_To_Sram_FIFO_18[15];
        Psram_En_To_Sram_FIFO_19[14] <= Psram_En_To_Sram_FIFO_19[15];
        Psram_En_To_Sram_FIFO_20[14] <= Psram_En_To_Sram_FIFO_20[15];
        Psram_En_To_Sram_FIFO_21[14] <= Psram_En_To_Sram_FIFO_21[15];
        Psram_En_To_Sram_FIFO_22[14] <= Psram_En_To_Sram_FIFO_22[15];
        Psram_En_To_Sram_FIFO_23[14] <= Psram_En_To_Sram_FIFO_23[15];
        Psram_En_To_Sram_FIFO_24[14] <= Psram_En_To_Sram_FIFO_24[15];
        Psram_En_To_Sram_FIFO_25[14] <= Psram_En_To_Sram_FIFO_25[15];
        Psram_En_To_Sram_FIFO_26[14] <= Psram_En_To_Sram_FIFO_26[15];
        Psram_En_To_Sram_FIFO_27[14] <= Psram_En_To_Sram_FIFO_27[15];
        Psram_En_To_Sram_FIFO_28[14] <= Psram_En_To_Sram_FIFO_28[15];
        Psram_En_To_Sram_FIFO_29[14] <= Psram_En_To_Sram_FIFO_29[15];
        Psram_En_To_Sram_FIFO_30[14] <= Psram_En_To_Sram_FIFO_30[15];
        Psram_En_To_Sram_FIFO_31[14] <= Psram_En_To_Sram_FIFO_31[15];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_16[15] <= i_Psram_En[16];
        Psram_En_To_Sram_FIFO_17[15] <= Psram_En_To_Sram_FIFO_17[16];
        Psram_En_To_Sram_FIFO_18[15] <= Psram_En_To_Sram_FIFO_18[16];
        Psram_En_To_Sram_FIFO_19[15] <= Psram_En_To_Sram_FIFO_19[16];
        Psram_En_To_Sram_FIFO_20[15] <= Psram_En_To_Sram_FIFO_20[16];
        Psram_En_To_Sram_FIFO_21[15] <= Psram_En_To_Sram_FIFO_21[16];
        Psram_En_To_Sram_FIFO_22[15] <= Psram_En_To_Sram_FIFO_22[16];
        Psram_En_To_Sram_FIFO_23[15] <= Psram_En_To_Sram_FIFO_23[16];
        Psram_En_To_Sram_FIFO_24[15] <= Psram_En_To_Sram_FIFO_24[16];
        Psram_En_To_Sram_FIFO_25[15] <= Psram_En_To_Sram_FIFO_25[16];
        Psram_En_To_Sram_FIFO_26[15] <= Psram_En_To_Sram_FIFO_26[16];
        Psram_En_To_Sram_FIFO_27[15] <= Psram_En_To_Sram_FIFO_27[16];
        Psram_En_To_Sram_FIFO_28[15] <= Psram_En_To_Sram_FIFO_28[16];
        Psram_En_To_Sram_FIFO_29[15] <= Psram_En_To_Sram_FIFO_29[16];
        Psram_En_To_Sram_FIFO_30[15] <= Psram_En_To_Sram_FIFO_30[16];
        Psram_En_To_Sram_FIFO_31[15] <= Psram_En_To_Sram_FIFO_31[16];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_17[16] <= i_Psram_En[17];
        Psram_En_To_Sram_FIFO_18[16] <= Psram_En_To_Sram_FIFO_18[17];
        Psram_En_To_Sram_FIFO_19[16] <= Psram_En_To_Sram_FIFO_19[17];
        Psram_En_To_Sram_FIFO_20[16] <= Psram_En_To_Sram_FIFO_20[17];
        Psram_En_To_Sram_FIFO_21[16] <= Psram_En_To_Sram_FIFO_21[17];
        Psram_En_To_Sram_FIFO_22[16] <= Psram_En_To_Sram_FIFO_22[17];
        Psram_En_To_Sram_FIFO_23[16] <= Psram_En_To_Sram_FIFO_23[17];
        Psram_En_To_Sram_FIFO_24[16] <= Psram_En_To_Sram_FIFO_24[17];
        Psram_En_To_Sram_FIFO_25[16] <= Psram_En_To_Sram_FIFO_25[17];
        Psram_En_To_Sram_FIFO_26[16] <= Psram_En_To_Sram_FIFO_26[17];
        Psram_En_To_Sram_FIFO_27[16] <= Psram_En_To_Sram_FIFO_27[17];
        Psram_En_To_Sram_FIFO_28[16] <= Psram_En_To_Sram_FIFO_28[17];
        Psram_En_To_Sram_FIFO_29[16] <= Psram_En_To_Sram_FIFO_29[17];
        Psram_En_To_Sram_FIFO_30[16] <= Psram_En_To_Sram_FIFO_30[17];
        Psram_En_To_Sram_FIFO_31[16] <= Psram_En_To_Sram_FIFO_31[17];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_18[17] <= i_Psram_En[18];
        Psram_En_To_Sram_FIFO_19[17] <= Psram_En_To_Sram_FIFO_19[18];
        Psram_En_To_Sram_FIFO_20[17] <= Psram_En_To_Sram_FIFO_20[18];
        Psram_En_To_Sram_FIFO_21[17] <= Psram_En_To_Sram_FIFO_21[18];
        Psram_En_To_Sram_FIFO_22[17] <= Psram_En_To_Sram_FIFO_22[18];
        Psram_En_To_Sram_FIFO_23[17] <= Psram_En_To_Sram_FIFO_23[18];
        Psram_En_To_Sram_FIFO_24[17] <= Psram_En_To_Sram_FIFO_24[18];
        Psram_En_To_Sram_FIFO_25[17] <= Psram_En_To_Sram_FIFO_25[18];
        Psram_En_To_Sram_FIFO_26[17] <= Psram_En_To_Sram_FIFO_26[18];
        Psram_En_To_Sram_FIFO_27[17] <= Psram_En_To_Sram_FIFO_27[18];
        Psram_En_To_Sram_FIFO_28[17] <= Psram_En_To_Sram_FIFO_28[18];
        Psram_En_To_Sram_FIFO_29[17] <= Psram_En_To_Sram_FIFO_29[18];
        Psram_En_To_Sram_FIFO_30[17] <= Psram_En_To_Sram_FIFO_30[18];
        Psram_En_To_Sram_FIFO_31[17] <= Psram_En_To_Sram_FIFO_31[18];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_19[18] <= i_Psram_En[19];
        Psram_En_To_Sram_FIFO_20[18] <= Psram_En_To_Sram_FIFO_20[19];
        Psram_En_To_Sram_FIFO_21[18] <= Psram_En_To_Sram_FIFO_21[19];
        Psram_En_To_Sram_FIFO_22[18] <= Psram_En_To_Sram_FIFO_22[19];
        Psram_En_To_Sram_FIFO_23[18] <= Psram_En_To_Sram_FIFO_23[19];
        Psram_En_To_Sram_FIFO_24[18] <= Psram_En_To_Sram_FIFO_24[19];
        Psram_En_To_Sram_FIFO_25[18] <= Psram_En_To_Sram_FIFO_25[19];
        Psram_En_To_Sram_FIFO_26[18] <= Psram_En_To_Sram_FIFO_26[19];
        Psram_En_To_Sram_FIFO_27[18] <= Psram_En_To_Sram_FIFO_27[19];
        Psram_En_To_Sram_FIFO_28[18] <= Psram_En_To_Sram_FIFO_28[19];
        Psram_En_To_Sram_FIFO_29[18] <= Psram_En_To_Sram_FIFO_29[19];
        Psram_En_To_Sram_FIFO_30[18] <= Psram_En_To_Sram_FIFO_30[19];
        Psram_En_To_Sram_FIFO_31[18] <= Psram_En_To_Sram_FIFO_31[19];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_20[19] <= i_Psram_En[20];
        Psram_En_To_Sram_FIFO_21[19] <= Psram_En_To_Sram_FIFO_21[20];
        Psram_En_To_Sram_FIFO_22[19] <= Psram_En_To_Sram_FIFO_22[20];
        Psram_En_To_Sram_FIFO_23[19] <= Psram_En_To_Sram_FIFO_23[20];
        Psram_En_To_Sram_FIFO_24[19] <= Psram_En_To_Sram_FIFO_24[20];
        Psram_En_To_Sram_FIFO_25[19] <= Psram_En_To_Sram_FIFO_25[20];
        Psram_En_To_Sram_FIFO_26[19] <= Psram_En_To_Sram_FIFO_26[20];
        Psram_En_To_Sram_FIFO_27[19] <= Psram_En_To_Sram_FIFO_27[20];
        Psram_En_To_Sram_FIFO_28[19] <= Psram_En_To_Sram_FIFO_28[20];
        Psram_En_To_Sram_FIFO_29[19] <= Psram_En_To_Sram_FIFO_29[20];
        Psram_En_To_Sram_FIFO_30[19] <= Psram_En_To_Sram_FIFO_30[20];
        Psram_En_To_Sram_FIFO_31[19] <= Psram_En_To_Sram_FIFO_31[20];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_21[20] <= i_Psram_En[21];
        Psram_En_To_Sram_FIFO_22[20] <= Psram_En_To_Sram_FIFO_22[21];
        Psram_En_To_Sram_FIFO_23[20] <= Psram_En_To_Sram_FIFO_23[21];
        Psram_En_To_Sram_FIFO_24[20] <= Psram_En_To_Sram_FIFO_24[21];
        Psram_En_To_Sram_FIFO_25[20] <= Psram_En_To_Sram_FIFO_25[21];
        Psram_En_To_Sram_FIFO_26[20] <= Psram_En_To_Sram_FIFO_26[21];
        Psram_En_To_Sram_FIFO_27[20] <= Psram_En_To_Sram_FIFO_27[21];
        Psram_En_To_Sram_FIFO_28[20] <= Psram_En_To_Sram_FIFO_28[21];
        Psram_En_To_Sram_FIFO_29[20] <= Psram_En_To_Sram_FIFO_29[21];
        Psram_En_To_Sram_FIFO_30[20] <= Psram_En_To_Sram_FIFO_30[21];
        Psram_En_To_Sram_FIFO_31[20] <= Psram_En_To_Sram_FIFO_31[21];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_22[21] <= i_Psram_En[22];
        Psram_En_To_Sram_FIFO_23[21] <= Psram_En_To_Sram_FIFO_23[22];
        Psram_En_To_Sram_FIFO_24[21] <= Psram_En_To_Sram_FIFO_24[22];
        Psram_En_To_Sram_FIFO_25[21] <= Psram_En_To_Sram_FIFO_25[22];
        Psram_En_To_Sram_FIFO_26[21] <= Psram_En_To_Sram_FIFO_26[22];
        Psram_En_To_Sram_FIFO_27[21] <= Psram_En_To_Sram_FIFO_27[22];
        Psram_En_To_Sram_FIFO_28[21] <= Psram_En_To_Sram_FIFO_28[22];
        Psram_En_To_Sram_FIFO_29[21] <= Psram_En_To_Sram_FIFO_29[22];
        Psram_En_To_Sram_FIFO_30[21] <= Psram_En_To_Sram_FIFO_30[22];
        Psram_En_To_Sram_FIFO_31[21] <= Psram_En_To_Sram_FIFO_31[22];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_23[22] <= i_Psram_En[23];
        Psram_En_To_Sram_FIFO_24[22] <= Psram_En_To_Sram_FIFO_24[23];
        Psram_En_To_Sram_FIFO_25[22] <= Psram_En_To_Sram_FIFO_25[23];
        Psram_En_To_Sram_FIFO_26[22] <= Psram_En_To_Sram_FIFO_26[23];
        Psram_En_To_Sram_FIFO_27[22] <= Psram_En_To_Sram_FIFO_27[23];
        Psram_En_To_Sram_FIFO_28[22] <= Psram_En_To_Sram_FIFO_28[23];
        Psram_En_To_Sram_FIFO_29[22] <= Psram_En_To_Sram_FIFO_29[23];
        Psram_En_To_Sram_FIFO_30[22] <= Psram_En_To_Sram_FIFO_30[23];
        Psram_En_To_Sram_FIFO_31[22] <= Psram_En_To_Sram_FIFO_31[23];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_24[23] <= i_Psram_En[24];
        Psram_En_To_Sram_FIFO_25[23] <= Psram_En_To_Sram_FIFO_25[24];
        Psram_En_To_Sram_FIFO_26[23] <= Psram_En_To_Sram_FIFO_26[24];
        Psram_En_To_Sram_FIFO_27[23] <= Psram_En_To_Sram_FIFO_27[24];
        Psram_En_To_Sram_FIFO_28[23] <= Psram_En_To_Sram_FIFO_28[24];
        Psram_En_To_Sram_FIFO_29[23] <= Psram_En_To_Sram_FIFO_29[24];
        Psram_En_To_Sram_FIFO_30[23] <= Psram_En_To_Sram_FIFO_30[24];
        Psram_En_To_Sram_FIFO_31[23] <= Psram_En_To_Sram_FIFO_31[24];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_25[24] <= i_Psram_En[25];
        Psram_En_To_Sram_FIFO_26[24] <= Psram_En_To_Sram_FIFO_26[25];
        Psram_En_To_Sram_FIFO_27[24] <= Psram_En_To_Sram_FIFO_27[25];
        Psram_En_To_Sram_FIFO_28[24] <= Psram_En_To_Sram_FIFO_28[25];
        Psram_En_To_Sram_FIFO_29[24] <= Psram_En_To_Sram_FIFO_29[25];
        Psram_En_To_Sram_FIFO_30[24] <= Psram_En_To_Sram_FIFO_30[25];
        Psram_En_To_Sram_FIFO_31[24] <= Psram_En_To_Sram_FIFO_31[25];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_26[25] <= i_Psram_En[26];
        Psram_En_To_Sram_FIFO_27[25] <= Psram_En_To_Sram_FIFO_27[26];
        Psram_En_To_Sram_FIFO_28[25] <= Psram_En_To_Sram_FIFO_28[26];
        Psram_En_To_Sram_FIFO_29[25] <= Psram_En_To_Sram_FIFO_29[26];
        Psram_En_To_Sram_FIFO_30[25] <= Psram_En_To_Sram_FIFO_30[26];
        Psram_En_To_Sram_FIFO_31[25] <= Psram_En_To_Sram_FIFO_31[26];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_27[26] <= i_Psram_En[27];
        Psram_En_To_Sram_FIFO_28[26] <= Psram_En_To_Sram_FIFO_28[27];
        Psram_En_To_Sram_FIFO_29[26] <= Psram_En_To_Sram_FIFO_29[27];
        Psram_En_To_Sram_FIFO_30[26] <= Psram_En_To_Sram_FIFO_30[27];
        Psram_En_To_Sram_FIFO_31[26] <= Psram_En_To_Sram_FIFO_31[27];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_28[27] <= i_Psram_En[28];
        Psram_En_To_Sram_FIFO_29[27] <= Psram_En_To_Sram_FIFO_29[28];
        Psram_En_To_Sram_FIFO_30[27] <= Psram_En_To_Sram_FIFO_30[28];
        Psram_En_To_Sram_FIFO_31[27] <= Psram_En_To_Sram_FIFO_31[28];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_29[28] <= i_Psram_En[29];
        Psram_En_To_Sram_FIFO_30[28] <= Psram_En_To_Sram_FIFO_30[29];
        Psram_En_To_Sram_FIFO_31[28] <= Psram_En_To_Sram_FIFO_31[29];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_30[29] <= i_Psram_En[30];
        Psram_En_To_Sram_FIFO_31[29] <= Psram_En_To_Sram_FIFO_31[30];
    end

    always @(posedge CLK) begin
        Psram_En_To_Sram_FIFO_31[30] <= i_Psram_En[31];
    end

    // Psram_Valid_To_Systolic Logic
    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_1[0] <= i_Psram_Valid_1buf[1];
        Psram_Valid_To_Systolic_FIFO_2[0] <= Psram_Valid_To_Systolic_FIFO_2[1];
        Psram_Valid_To_Systolic_FIFO_3[0] <= Psram_Valid_To_Systolic_FIFO_3[1];
        Psram_Valid_To_Systolic_FIFO_4[0] <= Psram_Valid_To_Systolic_FIFO_4[1];
        Psram_Valid_To_Systolic_FIFO_5[0] <= Psram_Valid_To_Systolic_FIFO_5[1];
        Psram_Valid_To_Systolic_FIFO_6[0] <= Psram_Valid_To_Systolic_FIFO_6[1];
        Psram_Valid_To_Systolic_FIFO_7[0] <= Psram_Valid_To_Systolic_FIFO_7[1];
        Psram_Valid_To_Systolic_FIFO_8[0] <= Psram_Valid_To_Systolic_FIFO_8[1];
        Psram_Valid_To_Systolic_FIFO_9[0] <= Psram_Valid_To_Systolic_FIFO_9[1];
        Psram_Valid_To_Systolic_FIFO_10[0] <= Psram_Valid_To_Systolic_FIFO_10[1];
        Psram_Valid_To_Systolic_FIFO_11[0] <= Psram_Valid_To_Systolic_FIFO_11[1];
        Psram_Valid_To_Systolic_FIFO_12[0] <= Psram_Valid_To_Systolic_FIFO_12[1];
        Psram_Valid_To_Systolic_FIFO_13[0] <= Psram_Valid_To_Systolic_FIFO_13[1];
        Psram_Valid_To_Systolic_FIFO_14[0] <= Psram_Valid_To_Systolic_FIFO_14[1];
        Psram_Valid_To_Systolic_FIFO_15[0] <= Psram_Valid_To_Systolic_FIFO_15[1];
        Psram_Valid_To_Systolic_FIFO_16[0] <= Psram_Valid_To_Systolic_FIFO_16[1];
        Psram_Valid_To_Systolic_FIFO_17[0] <= Psram_Valid_To_Systolic_FIFO_17[1];
        Psram_Valid_To_Systolic_FIFO_18[0] <= Psram_Valid_To_Systolic_FIFO_18[1];
        Psram_Valid_To_Systolic_FIFO_19[0] <= Psram_Valid_To_Systolic_FIFO_19[1];
        Psram_Valid_To_Systolic_FIFO_20[0] <= Psram_Valid_To_Systolic_FIFO_20[1];
        Psram_Valid_To_Systolic_FIFO_21[0] <= Psram_Valid_To_Systolic_FIFO_21[1];
        Psram_Valid_To_Systolic_FIFO_22[0] <= Psram_Valid_To_Systolic_FIFO_22[1];
        Psram_Valid_To_Systolic_FIFO_23[0] <= Psram_Valid_To_Systolic_FIFO_23[1];
        Psram_Valid_To_Systolic_FIFO_24[0] <= Psram_Valid_To_Systolic_FIFO_24[1];
        Psram_Valid_To_Systolic_FIFO_25[0] <= Psram_Valid_To_Systolic_FIFO_25[1];
        Psram_Valid_To_Systolic_FIFO_26[0] <= Psram_Valid_To_Systolic_FIFO_26[1];
        Psram_Valid_To_Systolic_FIFO_27[0] <= Psram_Valid_To_Systolic_FIFO_27[1];
        Psram_Valid_To_Systolic_FIFO_28[0] <= Psram_Valid_To_Systolic_FIFO_28[1];
        Psram_Valid_To_Systolic_FIFO_29[0] <= Psram_Valid_To_Systolic_FIFO_29[1];
        Psram_Valid_To_Systolic_FIFO_30[0] <= Psram_Valid_To_Systolic_FIFO_30[1];
        Psram_Valid_To_Systolic_FIFO_31[0] <= Psram_Valid_To_Systolic_FIFO_31[1];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_2[1] <= i_Psram_Valid_1buf[2];
        Psram_Valid_To_Systolic_FIFO_3[1] <= Psram_Valid_To_Systolic_FIFO_3[2];
        Psram_Valid_To_Systolic_FIFO_4[1] <= Psram_Valid_To_Systolic_FIFO_4[2];
        Psram_Valid_To_Systolic_FIFO_5[1] <= Psram_Valid_To_Systolic_FIFO_5[2];
        Psram_Valid_To_Systolic_FIFO_6[1] <= Psram_Valid_To_Systolic_FIFO_6[2];
        Psram_Valid_To_Systolic_FIFO_7[1] <= Psram_Valid_To_Systolic_FIFO_7[2];
        Psram_Valid_To_Systolic_FIFO_8[1] <= Psram_Valid_To_Systolic_FIFO_8[2];
        Psram_Valid_To_Systolic_FIFO_9[1] <= Psram_Valid_To_Systolic_FIFO_9[2];
        Psram_Valid_To_Systolic_FIFO_10[1] <= Psram_Valid_To_Systolic_FIFO_10[2];
        Psram_Valid_To_Systolic_FIFO_11[1] <= Psram_Valid_To_Systolic_FIFO_11[2];
        Psram_Valid_To_Systolic_FIFO_12[1] <= Psram_Valid_To_Systolic_FIFO_12[2];
        Psram_Valid_To_Systolic_FIFO_13[1] <= Psram_Valid_To_Systolic_FIFO_13[2];
        Psram_Valid_To_Systolic_FIFO_14[1] <= Psram_Valid_To_Systolic_FIFO_14[2];
        Psram_Valid_To_Systolic_FIFO_15[1] <= Psram_Valid_To_Systolic_FIFO_15[2];
        Psram_Valid_To_Systolic_FIFO_16[1] <= Psram_Valid_To_Systolic_FIFO_16[2];
        Psram_Valid_To_Systolic_FIFO_17[1] <= Psram_Valid_To_Systolic_FIFO_17[2];
        Psram_Valid_To_Systolic_FIFO_18[1] <= Psram_Valid_To_Systolic_FIFO_18[2];
        Psram_Valid_To_Systolic_FIFO_19[1] <= Psram_Valid_To_Systolic_FIFO_19[2];
        Psram_Valid_To_Systolic_FIFO_20[1] <= Psram_Valid_To_Systolic_FIFO_20[2];
        Psram_Valid_To_Systolic_FIFO_21[1] <= Psram_Valid_To_Systolic_FIFO_21[2];
        Psram_Valid_To_Systolic_FIFO_22[1] <= Psram_Valid_To_Systolic_FIFO_22[2];
        Psram_Valid_To_Systolic_FIFO_23[1] <= Psram_Valid_To_Systolic_FIFO_23[2];
        Psram_Valid_To_Systolic_FIFO_24[1] <= Psram_Valid_To_Systolic_FIFO_24[2];
        Psram_Valid_To_Systolic_FIFO_25[1] <= Psram_Valid_To_Systolic_FIFO_25[2];
        Psram_Valid_To_Systolic_FIFO_26[1] <= Psram_Valid_To_Systolic_FIFO_26[2];
        Psram_Valid_To_Systolic_FIFO_27[1] <= Psram_Valid_To_Systolic_FIFO_27[2];
        Psram_Valid_To_Systolic_FIFO_28[1] <= Psram_Valid_To_Systolic_FIFO_28[2];
        Psram_Valid_To_Systolic_FIFO_29[1] <= Psram_Valid_To_Systolic_FIFO_29[2];
        Psram_Valid_To_Systolic_FIFO_30[1] <= Psram_Valid_To_Systolic_FIFO_30[2];
        Psram_Valid_To_Systolic_FIFO_31[1] <= Psram_Valid_To_Systolic_FIFO_31[2];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_3[2] <= i_Psram_Valid_1buf[3];
        Psram_Valid_To_Systolic_FIFO_4[2] <= Psram_Valid_To_Systolic_FIFO_4[3];
        Psram_Valid_To_Systolic_FIFO_5[2] <= Psram_Valid_To_Systolic_FIFO_5[3];
        Psram_Valid_To_Systolic_FIFO_6[2] <= Psram_Valid_To_Systolic_FIFO_6[3];
        Psram_Valid_To_Systolic_FIFO_7[2] <= Psram_Valid_To_Systolic_FIFO_7[3];
        Psram_Valid_To_Systolic_FIFO_8[2] <= Psram_Valid_To_Systolic_FIFO_8[3];
        Psram_Valid_To_Systolic_FIFO_9[2] <= Psram_Valid_To_Systolic_FIFO_9[3];
        Psram_Valid_To_Systolic_FIFO_10[2] <= Psram_Valid_To_Systolic_FIFO_10[3];
        Psram_Valid_To_Systolic_FIFO_11[2] <= Psram_Valid_To_Systolic_FIFO_11[3];
        Psram_Valid_To_Systolic_FIFO_12[2] <= Psram_Valid_To_Systolic_FIFO_12[3];
        Psram_Valid_To_Systolic_FIFO_13[2] <= Psram_Valid_To_Systolic_FIFO_13[3];
        Psram_Valid_To_Systolic_FIFO_14[2] <= Psram_Valid_To_Systolic_FIFO_14[3];
        Psram_Valid_To_Systolic_FIFO_15[2] <= Psram_Valid_To_Systolic_FIFO_15[3];
        Psram_Valid_To_Systolic_FIFO_16[2] <= Psram_Valid_To_Systolic_FIFO_16[3];
        Psram_Valid_To_Systolic_FIFO_17[2] <= Psram_Valid_To_Systolic_FIFO_17[3];
        Psram_Valid_To_Systolic_FIFO_18[2] <= Psram_Valid_To_Systolic_FIFO_18[3];
        Psram_Valid_To_Systolic_FIFO_19[2] <= Psram_Valid_To_Systolic_FIFO_19[3];
        Psram_Valid_To_Systolic_FIFO_20[2] <= Psram_Valid_To_Systolic_FIFO_20[3];
        Psram_Valid_To_Systolic_FIFO_21[2] <= Psram_Valid_To_Systolic_FIFO_21[3];
        Psram_Valid_To_Systolic_FIFO_22[2] <= Psram_Valid_To_Systolic_FIFO_22[3];
        Psram_Valid_To_Systolic_FIFO_23[2] <= Psram_Valid_To_Systolic_FIFO_23[3];
        Psram_Valid_To_Systolic_FIFO_24[2] <= Psram_Valid_To_Systolic_FIFO_24[3];
        Psram_Valid_To_Systolic_FIFO_25[2] <= Psram_Valid_To_Systolic_FIFO_25[3];
        Psram_Valid_To_Systolic_FIFO_26[2] <= Psram_Valid_To_Systolic_FIFO_26[3];
        Psram_Valid_To_Systolic_FIFO_27[2] <= Psram_Valid_To_Systolic_FIFO_27[3];
        Psram_Valid_To_Systolic_FIFO_28[2] <= Psram_Valid_To_Systolic_FIFO_28[3];
        Psram_Valid_To_Systolic_FIFO_29[2] <= Psram_Valid_To_Systolic_FIFO_29[3];
        Psram_Valid_To_Systolic_FIFO_30[2] <= Psram_Valid_To_Systolic_FIFO_30[3];
        Psram_Valid_To_Systolic_FIFO_31[2] <= Psram_Valid_To_Systolic_FIFO_31[3];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_4[3] <= i_Psram_Valid_1buf[4];
        Psram_Valid_To_Systolic_FIFO_5[3] <= Psram_Valid_To_Systolic_FIFO_5[4];
        Psram_Valid_To_Systolic_FIFO_6[3] <= Psram_Valid_To_Systolic_FIFO_6[4];
        Psram_Valid_To_Systolic_FIFO_7[3] <= Psram_Valid_To_Systolic_FIFO_7[4];
        Psram_Valid_To_Systolic_FIFO_8[3] <= Psram_Valid_To_Systolic_FIFO_8[4];
        Psram_Valid_To_Systolic_FIFO_9[3] <= Psram_Valid_To_Systolic_FIFO_9[4];
        Psram_Valid_To_Systolic_FIFO_10[3] <= Psram_Valid_To_Systolic_FIFO_10[4];
        Psram_Valid_To_Systolic_FIFO_11[3] <= Psram_Valid_To_Systolic_FIFO_11[4];
        Psram_Valid_To_Systolic_FIFO_12[3] <= Psram_Valid_To_Systolic_FIFO_12[4];
        Psram_Valid_To_Systolic_FIFO_13[3] <= Psram_Valid_To_Systolic_FIFO_13[4];
        Psram_Valid_To_Systolic_FIFO_14[3] <= Psram_Valid_To_Systolic_FIFO_14[4];
        Psram_Valid_To_Systolic_FIFO_15[3] <= Psram_Valid_To_Systolic_FIFO_15[4];
        Psram_Valid_To_Systolic_FIFO_16[3] <= Psram_Valid_To_Systolic_FIFO_16[4];
        Psram_Valid_To_Systolic_FIFO_17[3] <= Psram_Valid_To_Systolic_FIFO_17[4];
        Psram_Valid_To_Systolic_FIFO_18[3] <= Psram_Valid_To_Systolic_FIFO_18[4];
        Psram_Valid_To_Systolic_FIFO_19[3] <= Psram_Valid_To_Systolic_FIFO_19[4];
        Psram_Valid_To_Systolic_FIFO_20[3] <= Psram_Valid_To_Systolic_FIFO_20[4];
        Psram_Valid_To_Systolic_FIFO_21[3] <= Psram_Valid_To_Systolic_FIFO_21[4];
        Psram_Valid_To_Systolic_FIFO_22[3] <= Psram_Valid_To_Systolic_FIFO_22[4];
        Psram_Valid_To_Systolic_FIFO_23[3] <= Psram_Valid_To_Systolic_FIFO_23[4];
        Psram_Valid_To_Systolic_FIFO_24[3] <= Psram_Valid_To_Systolic_FIFO_24[4];
        Psram_Valid_To_Systolic_FIFO_25[3] <= Psram_Valid_To_Systolic_FIFO_25[4];
        Psram_Valid_To_Systolic_FIFO_26[3] <= Psram_Valid_To_Systolic_FIFO_26[4];
        Psram_Valid_To_Systolic_FIFO_27[3] <= Psram_Valid_To_Systolic_FIFO_27[4];
        Psram_Valid_To_Systolic_FIFO_28[3] <= Psram_Valid_To_Systolic_FIFO_28[4];
        Psram_Valid_To_Systolic_FIFO_29[3] <= Psram_Valid_To_Systolic_FIFO_29[4];
        Psram_Valid_To_Systolic_FIFO_30[3] <= Psram_Valid_To_Systolic_FIFO_30[4];
        Psram_Valid_To_Systolic_FIFO_31[3] <= Psram_Valid_To_Systolic_FIFO_31[4];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_5[4] <= i_Psram_Valid_1buf[5];
        Psram_Valid_To_Systolic_FIFO_6[4] <= Psram_Valid_To_Systolic_FIFO_6[5];
        Psram_Valid_To_Systolic_FIFO_7[4] <= Psram_Valid_To_Systolic_FIFO_7[5];
        Psram_Valid_To_Systolic_FIFO_8[4] <= Psram_Valid_To_Systolic_FIFO_8[5];
        Psram_Valid_To_Systolic_FIFO_9[4] <= Psram_Valid_To_Systolic_FIFO_9[5];
        Psram_Valid_To_Systolic_FIFO_10[4] <= Psram_Valid_To_Systolic_FIFO_10[5];
        Psram_Valid_To_Systolic_FIFO_11[4] <= Psram_Valid_To_Systolic_FIFO_11[5];
        Psram_Valid_To_Systolic_FIFO_12[4] <= Psram_Valid_To_Systolic_FIFO_12[5];
        Psram_Valid_To_Systolic_FIFO_13[4] <= Psram_Valid_To_Systolic_FIFO_13[5];
        Psram_Valid_To_Systolic_FIFO_14[4] <= Psram_Valid_To_Systolic_FIFO_14[5];
        Psram_Valid_To_Systolic_FIFO_15[4] <= Psram_Valid_To_Systolic_FIFO_15[5];
        Psram_Valid_To_Systolic_FIFO_16[4] <= Psram_Valid_To_Systolic_FIFO_16[5];
        Psram_Valid_To_Systolic_FIFO_17[4] <= Psram_Valid_To_Systolic_FIFO_17[5];
        Psram_Valid_To_Systolic_FIFO_18[4] <= Psram_Valid_To_Systolic_FIFO_18[5];
        Psram_Valid_To_Systolic_FIFO_19[4] <= Psram_Valid_To_Systolic_FIFO_19[5];
        Psram_Valid_To_Systolic_FIFO_20[4] <= Psram_Valid_To_Systolic_FIFO_20[5];
        Psram_Valid_To_Systolic_FIFO_21[4] <= Psram_Valid_To_Systolic_FIFO_21[5];
        Psram_Valid_To_Systolic_FIFO_22[4] <= Psram_Valid_To_Systolic_FIFO_22[5];
        Psram_Valid_To_Systolic_FIFO_23[4] <= Psram_Valid_To_Systolic_FIFO_23[5];
        Psram_Valid_To_Systolic_FIFO_24[4] <= Psram_Valid_To_Systolic_FIFO_24[5];
        Psram_Valid_To_Systolic_FIFO_25[4] <= Psram_Valid_To_Systolic_FIFO_25[5];
        Psram_Valid_To_Systolic_FIFO_26[4] <= Psram_Valid_To_Systolic_FIFO_26[5];
        Psram_Valid_To_Systolic_FIFO_27[4] <= Psram_Valid_To_Systolic_FIFO_27[5];
        Psram_Valid_To_Systolic_FIFO_28[4] <= Psram_Valid_To_Systolic_FIFO_28[5];
        Psram_Valid_To_Systolic_FIFO_29[4] <= Psram_Valid_To_Systolic_FIFO_29[5];
        Psram_Valid_To_Systolic_FIFO_30[4] <= Psram_Valid_To_Systolic_FIFO_30[5];
        Psram_Valid_To_Systolic_FIFO_31[4] <= Psram_Valid_To_Systolic_FIFO_31[5];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_6[5] <= i_Psram_Valid_1buf[6];
        Psram_Valid_To_Systolic_FIFO_7[5] <= Psram_Valid_To_Systolic_FIFO_7[6];
        Psram_Valid_To_Systolic_FIFO_8[5] <= Psram_Valid_To_Systolic_FIFO_8[6];
        Psram_Valid_To_Systolic_FIFO_9[5] <= Psram_Valid_To_Systolic_FIFO_9[6];
        Psram_Valid_To_Systolic_FIFO_10[5] <= Psram_Valid_To_Systolic_FIFO_10[6];
        Psram_Valid_To_Systolic_FIFO_11[5] <= Psram_Valid_To_Systolic_FIFO_11[6];
        Psram_Valid_To_Systolic_FIFO_12[5] <= Psram_Valid_To_Systolic_FIFO_12[6];
        Psram_Valid_To_Systolic_FIFO_13[5] <= Psram_Valid_To_Systolic_FIFO_13[6];
        Psram_Valid_To_Systolic_FIFO_14[5] <= Psram_Valid_To_Systolic_FIFO_14[6];
        Psram_Valid_To_Systolic_FIFO_15[5] <= Psram_Valid_To_Systolic_FIFO_15[6];
        Psram_Valid_To_Systolic_FIFO_16[5] <= Psram_Valid_To_Systolic_FIFO_16[6];
        Psram_Valid_To_Systolic_FIFO_17[5] <= Psram_Valid_To_Systolic_FIFO_17[6];
        Psram_Valid_To_Systolic_FIFO_18[5] <= Psram_Valid_To_Systolic_FIFO_18[6];
        Psram_Valid_To_Systolic_FIFO_19[5] <= Psram_Valid_To_Systolic_FIFO_19[6];
        Psram_Valid_To_Systolic_FIFO_20[5] <= Psram_Valid_To_Systolic_FIFO_20[6];
        Psram_Valid_To_Systolic_FIFO_21[5] <= Psram_Valid_To_Systolic_FIFO_21[6];
        Psram_Valid_To_Systolic_FIFO_22[5] <= Psram_Valid_To_Systolic_FIFO_22[6];
        Psram_Valid_To_Systolic_FIFO_23[5] <= Psram_Valid_To_Systolic_FIFO_23[6];
        Psram_Valid_To_Systolic_FIFO_24[5] <= Psram_Valid_To_Systolic_FIFO_24[6];
        Psram_Valid_To_Systolic_FIFO_25[5] <= Psram_Valid_To_Systolic_FIFO_25[6];
        Psram_Valid_To_Systolic_FIFO_26[5] <= Psram_Valid_To_Systolic_FIFO_26[6];
        Psram_Valid_To_Systolic_FIFO_27[5] <= Psram_Valid_To_Systolic_FIFO_27[6];
        Psram_Valid_To_Systolic_FIFO_28[5] <= Psram_Valid_To_Systolic_FIFO_28[6];
        Psram_Valid_To_Systolic_FIFO_29[5] <= Psram_Valid_To_Systolic_FIFO_29[6];
        Psram_Valid_To_Systolic_FIFO_30[5] <= Psram_Valid_To_Systolic_FIFO_30[6];
        Psram_Valid_To_Systolic_FIFO_31[5] <= Psram_Valid_To_Systolic_FIFO_31[6];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_7[6] <= i_Psram_Valid_1buf[7];
        Psram_Valid_To_Systolic_FIFO_8[6] <= Psram_Valid_To_Systolic_FIFO_8[7];
        Psram_Valid_To_Systolic_FIFO_9[6] <= Psram_Valid_To_Systolic_FIFO_9[7];
        Psram_Valid_To_Systolic_FIFO_10[6] <= Psram_Valid_To_Systolic_FIFO_10[7];
        Psram_Valid_To_Systolic_FIFO_11[6] <= Psram_Valid_To_Systolic_FIFO_11[7];
        Psram_Valid_To_Systolic_FIFO_12[6] <= Psram_Valid_To_Systolic_FIFO_12[7];
        Psram_Valid_To_Systolic_FIFO_13[6] <= Psram_Valid_To_Systolic_FIFO_13[7];
        Psram_Valid_To_Systolic_FIFO_14[6] <= Psram_Valid_To_Systolic_FIFO_14[7];
        Psram_Valid_To_Systolic_FIFO_15[6] <= Psram_Valid_To_Systolic_FIFO_15[7];
        Psram_Valid_To_Systolic_FIFO_16[6] <= Psram_Valid_To_Systolic_FIFO_16[7];
        Psram_Valid_To_Systolic_FIFO_17[6] <= Psram_Valid_To_Systolic_FIFO_17[7];
        Psram_Valid_To_Systolic_FIFO_18[6] <= Psram_Valid_To_Systolic_FIFO_18[7];
        Psram_Valid_To_Systolic_FIFO_19[6] <= Psram_Valid_To_Systolic_FIFO_19[7];
        Psram_Valid_To_Systolic_FIFO_20[6] <= Psram_Valid_To_Systolic_FIFO_20[7];
        Psram_Valid_To_Systolic_FIFO_21[6] <= Psram_Valid_To_Systolic_FIFO_21[7];
        Psram_Valid_To_Systolic_FIFO_22[6] <= Psram_Valid_To_Systolic_FIFO_22[7];
        Psram_Valid_To_Systolic_FIFO_23[6] <= Psram_Valid_To_Systolic_FIFO_23[7];
        Psram_Valid_To_Systolic_FIFO_24[6] <= Psram_Valid_To_Systolic_FIFO_24[7];
        Psram_Valid_To_Systolic_FIFO_25[6] <= Psram_Valid_To_Systolic_FIFO_25[7];
        Psram_Valid_To_Systolic_FIFO_26[6] <= Psram_Valid_To_Systolic_FIFO_26[7];
        Psram_Valid_To_Systolic_FIFO_27[6] <= Psram_Valid_To_Systolic_FIFO_27[7];
        Psram_Valid_To_Systolic_FIFO_28[6] <= Psram_Valid_To_Systolic_FIFO_28[7];
        Psram_Valid_To_Systolic_FIFO_29[6] <= Psram_Valid_To_Systolic_FIFO_29[7];
        Psram_Valid_To_Systolic_FIFO_30[6] <= Psram_Valid_To_Systolic_FIFO_30[7];
        Psram_Valid_To_Systolic_FIFO_31[6] <= Psram_Valid_To_Systolic_FIFO_31[7];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_8[7] <= i_Psram_Valid_1buf[8];
        Psram_Valid_To_Systolic_FIFO_9[7] <= Psram_Valid_To_Systolic_FIFO_9[8];
        Psram_Valid_To_Systolic_FIFO_10[7] <= Psram_Valid_To_Systolic_FIFO_10[8];
        Psram_Valid_To_Systolic_FIFO_11[7] <= Psram_Valid_To_Systolic_FIFO_11[8];
        Psram_Valid_To_Systolic_FIFO_12[7] <= Psram_Valid_To_Systolic_FIFO_12[8];
        Psram_Valid_To_Systolic_FIFO_13[7] <= Psram_Valid_To_Systolic_FIFO_13[8];
        Psram_Valid_To_Systolic_FIFO_14[7] <= Psram_Valid_To_Systolic_FIFO_14[8];
        Psram_Valid_To_Systolic_FIFO_15[7] <= Psram_Valid_To_Systolic_FIFO_15[8];
        Psram_Valid_To_Systolic_FIFO_16[7] <= Psram_Valid_To_Systolic_FIFO_16[8];
        Psram_Valid_To_Systolic_FIFO_17[7] <= Psram_Valid_To_Systolic_FIFO_17[8];
        Psram_Valid_To_Systolic_FIFO_18[7] <= Psram_Valid_To_Systolic_FIFO_18[8];
        Psram_Valid_To_Systolic_FIFO_19[7] <= Psram_Valid_To_Systolic_FIFO_19[8];
        Psram_Valid_To_Systolic_FIFO_20[7] <= Psram_Valid_To_Systolic_FIFO_20[8];
        Psram_Valid_To_Systolic_FIFO_21[7] <= Psram_Valid_To_Systolic_FIFO_21[8];
        Psram_Valid_To_Systolic_FIFO_22[7] <= Psram_Valid_To_Systolic_FIFO_22[8];
        Psram_Valid_To_Systolic_FIFO_23[7] <= Psram_Valid_To_Systolic_FIFO_23[8];
        Psram_Valid_To_Systolic_FIFO_24[7] <= Psram_Valid_To_Systolic_FIFO_24[8];
        Psram_Valid_To_Systolic_FIFO_25[7] <= Psram_Valid_To_Systolic_FIFO_25[8];
        Psram_Valid_To_Systolic_FIFO_26[7] <= Psram_Valid_To_Systolic_FIFO_26[8];
        Psram_Valid_To_Systolic_FIFO_27[7] <= Psram_Valid_To_Systolic_FIFO_27[8];
        Psram_Valid_To_Systolic_FIFO_28[7] <= Psram_Valid_To_Systolic_FIFO_28[8];
        Psram_Valid_To_Systolic_FIFO_29[7] <= Psram_Valid_To_Systolic_FIFO_29[8];
        Psram_Valid_To_Systolic_FIFO_30[7] <= Psram_Valid_To_Systolic_FIFO_30[8];
        Psram_Valid_To_Systolic_FIFO_31[7] <= Psram_Valid_To_Systolic_FIFO_31[8];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_9[8] <= i_Psram_Valid_1buf[9];
        Psram_Valid_To_Systolic_FIFO_10[8] <= Psram_Valid_To_Systolic_FIFO_10[9];
        Psram_Valid_To_Systolic_FIFO_11[8] <= Psram_Valid_To_Systolic_FIFO_11[9];
        Psram_Valid_To_Systolic_FIFO_12[8] <= Psram_Valid_To_Systolic_FIFO_12[9];
        Psram_Valid_To_Systolic_FIFO_13[8] <= Psram_Valid_To_Systolic_FIFO_13[9];
        Psram_Valid_To_Systolic_FIFO_14[8] <= Psram_Valid_To_Systolic_FIFO_14[9];
        Psram_Valid_To_Systolic_FIFO_15[8] <= Psram_Valid_To_Systolic_FIFO_15[9];
        Psram_Valid_To_Systolic_FIFO_16[8] <= Psram_Valid_To_Systolic_FIFO_16[9];
        Psram_Valid_To_Systolic_FIFO_17[8] <= Psram_Valid_To_Systolic_FIFO_17[9];
        Psram_Valid_To_Systolic_FIFO_18[8] <= Psram_Valid_To_Systolic_FIFO_18[9];
        Psram_Valid_To_Systolic_FIFO_19[8] <= Psram_Valid_To_Systolic_FIFO_19[9];
        Psram_Valid_To_Systolic_FIFO_20[8] <= Psram_Valid_To_Systolic_FIFO_20[9];
        Psram_Valid_To_Systolic_FIFO_21[8] <= Psram_Valid_To_Systolic_FIFO_21[9];
        Psram_Valid_To_Systolic_FIFO_22[8] <= Psram_Valid_To_Systolic_FIFO_22[9];
        Psram_Valid_To_Systolic_FIFO_23[8] <= Psram_Valid_To_Systolic_FIFO_23[9];
        Psram_Valid_To_Systolic_FIFO_24[8] <= Psram_Valid_To_Systolic_FIFO_24[9];
        Psram_Valid_To_Systolic_FIFO_25[8] <= Psram_Valid_To_Systolic_FIFO_25[9];
        Psram_Valid_To_Systolic_FIFO_26[8] <= Psram_Valid_To_Systolic_FIFO_26[9];
        Psram_Valid_To_Systolic_FIFO_27[8] <= Psram_Valid_To_Systolic_FIFO_27[9];
        Psram_Valid_To_Systolic_FIFO_28[8] <= Psram_Valid_To_Systolic_FIFO_28[9];
        Psram_Valid_To_Systolic_FIFO_29[8] <= Psram_Valid_To_Systolic_FIFO_29[9];
        Psram_Valid_To_Systolic_FIFO_30[8] <= Psram_Valid_To_Systolic_FIFO_30[9];
        Psram_Valid_To_Systolic_FIFO_31[8] <= Psram_Valid_To_Systolic_FIFO_31[9];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_10[9] <= i_Psram_Valid_1buf[10];
        Psram_Valid_To_Systolic_FIFO_11[9] <= Psram_Valid_To_Systolic_FIFO_11[10];
        Psram_Valid_To_Systolic_FIFO_12[9] <= Psram_Valid_To_Systolic_FIFO_12[10];
        Psram_Valid_To_Systolic_FIFO_13[9] <= Psram_Valid_To_Systolic_FIFO_13[10];
        Psram_Valid_To_Systolic_FIFO_14[9] <= Psram_Valid_To_Systolic_FIFO_14[10];
        Psram_Valid_To_Systolic_FIFO_15[9] <= Psram_Valid_To_Systolic_FIFO_15[10];
        Psram_Valid_To_Systolic_FIFO_16[9] <= Psram_Valid_To_Systolic_FIFO_16[10];
        Psram_Valid_To_Systolic_FIFO_17[9] <= Psram_Valid_To_Systolic_FIFO_17[10];
        Psram_Valid_To_Systolic_FIFO_18[9] <= Psram_Valid_To_Systolic_FIFO_18[10];
        Psram_Valid_To_Systolic_FIFO_19[9] <= Psram_Valid_To_Systolic_FIFO_19[10];
        Psram_Valid_To_Systolic_FIFO_20[9] <= Psram_Valid_To_Systolic_FIFO_20[10];
        Psram_Valid_To_Systolic_FIFO_21[9] <= Psram_Valid_To_Systolic_FIFO_21[10];
        Psram_Valid_To_Systolic_FIFO_22[9] <= Psram_Valid_To_Systolic_FIFO_22[10];
        Psram_Valid_To_Systolic_FIFO_23[9] <= Psram_Valid_To_Systolic_FIFO_23[10];
        Psram_Valid_To_Systolic_FIFO_24[9] <= Psram_Valid_To_Systolic_FIFO_24[10];
        Psram_Valid_To_Systolic_FIFO_25[9] <= Psram_Valid_To_Systolic_FIFO_25[10];
        Psram_Valid_To_Systolic_FIFO_26[9] <= Psram_Valid_To_Systolic_FIFO_26[10];
        Psram_Valid_To_Systolic_FIFO_27[9] <= Psram_Valid_To_Systolic_FIFO_27[10];
        Psram_Valid_To_Systolic_FIFO_28[9] <= Psram_Valid_To_Systolic_FIFO_28[10];
        Psram_Valid_To_Systolic_FIFO_29[9] <= Psram_Valid_To_Systolic_FIFO_29[10];
        Psram_Valid_To_Systolic_FIFO_30[9] <= Psram_Valid_To_Systolic_FIFO_30[10];
        Psram_Valid_To_Systolic_FIFO_31[9] <= Psram_Valid_To_Systolic_FIFO_31[10];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_11[10] <= i_Psram_Valid_1buf[11];
        Psram_Valid_To_Systolic_FIFO_12[10] <= Psram_Valid_To_Systolic_FIFO_12[11];
        Psram_Valid_To_Systolic_FIFO_13[10] <= Psram_Valid_To_Systolic_FIFO_13[11];
        Psram_Valid_To_Systolic_FIFO_14[10] <= Psram_Valid_To_Systolic_FIFO_14[11];
        Psram_Valid_To_Systolic_FIFO_15[10] <= Psram_Valid_To_Systolic_FIFO_15[11];
        Psram_Valid_To_Systolic_FIFO_16[10] <= Psram_Valid_To_Systolic_FIFO_16[11];
        Psram_Valid_To_Systolic_FIFO_17[10] <= Psram_Valid_To_Systolic_FIFO_17[11];
        Psram_Valid_To_Systolic_FIFO_18[10] <= Psram_Valid_To_Systolic_FIFO_18[11];
        Psram_Valid_To_Systolic_FIFO_19[10] <= Psram_Valid_To_Systolic_FIFO_19[11];
        Psram_Valid_To_Systolic_FIFO_20[10] <= Psram_Valid_To_Systolic_FIFO_20[11];
        Psram_Valid_To_Systolic_FIFO_21[10] <= Psram_Valid_To_Systolic_FIFO_21[11];
        Psram_Valid_To_Systolic_FIFO_22[10] <= Psram_Valid_To_Systolic_FIFO_22[11];
        Psram_Valid_To_Systolic_FIFO_23[10] <= Psram_Valid_To_Systolic_FIFO_23[11];
        Psram_Valid_To_Systolic_FIFO_24[10] <= Psram_Valid_To_Systolic_FIFO_24[11];
        Psram_Valid_To_Systolic_FIFO_25[10] <= Psram_Valid_To_Systolic_FIFO_25[11];
        Psram_Valid_To_Systolic_FIFO_26[10] <= Psram_Valid_To_Systolic_FIFO_26[11];
        Psram_Valid_To_Systolic_FIFO_27[10] <= Psram_Valid_To_Systolic_FIFO_27[11];
        Psram_Valid_To_Systolic_FIFO_28[10] <= Psram_Valid_To_Systolic_FIFO_28[11];
        Psram_Valid_To_Systolic_FIFO_29[10] <= Psram_Valid_To_Systolic_FIFO_29[11];
        Psram_Valid_To_Systolic_FIFO_30[10] <= Psram_Valid_To_Systolic_FIFO_30[11];
        Psram_Valid_To_Systolic_FIFO_31[10] <= Psram_Valid_To_Systolic_FIFO_31[11];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_12[11] <= i_Psram_Valid_1buf[12];
        Psram_Valid_To_Systolic_FIFO_13[11] <= Psram_Valid_To_Systolic_FIFO_13[12];
        Psram_Valid_To_Systolic_FIFO_14[11] <= Psram_Valid_To_Systolic_FIFO_14[12];
        Psram_Valid_To_Systolic_FIFO_15[11] <= Psram_Valid_To_Systolic_FIFO_15[12];
        Psram_Valid_To_Systolic_FIFO_16[11] <= Psram_Valid_To_Systolic_FIFO_16[12];
        Psram_Valid_To_Systolic_FIFO_17[11] <= Psram_Valid_To_Systolic_FIFO_17[12];
        Psram_Valid_To_Systolic_FIFO_18[11] <= Psram_Valid_To_Systolic_FIFO_18[12];
        Psram_Valid_To_Systolic_FIFO_19[11] <= Psram_Valid_To_Systolic_FIFO_19[12];
        Psram_Valid_To_Systolic_FIFO_20[11] <= Psram_Valid_To_Systolic_FIFO_20[12];
        Psram_Valid_To_Systolic_FIFO_21[11] <= Psram_Valid_To_Systolic_FIFO_21[12];
        Psram_Valid_To_Systolic_FIFO_22[11] <= Psram_Valid_To_Systolic_FIFO_22[12];
        Psram_Valid_To_Systolic_FIFO_23[11] <= Psram_Valid_To_Systolic_FIFO_23[12];
        Psram_Valid_To_Systolic_FIFO_24[11] <= Psram_Valid_To_Systolic_FIFO_24[12];
        Psram_Valid_To_Systolic_FIFO_25[11] <= Psram_Valid_To_Systolic_FIFO_25[12];
        Psram_Valid_To_Systolic_FIFO_26[11] <= Psram_Valid_To_Systolic_FIFO_26[12];
        Psram_Valid_To_Systolic_FIFO_27[11] <= Psram_Valid_To_Systolic_FIFO_27[12];
        Psram_Valid_To_Systolic_FIFO_28[11] <= Psram_Valid_To_Systolic_FIFO_28[12];
        Psram_Valid_To_Systolic_FIFO_29[11] <= Psram_Valid_To_Systolic_FIFO_29[12];
        Psram_Valid_To_Systolic_FIFO_30[11] <= Psram_Valid_To_Systolic_FIFO_30[12];
        Psram_Valid_To_Systolic_FIFO_31[11] <= Psram_Valid_To_Systolic_FIFO_31[12];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_13[12] <= i_Psram_Valid_1buf[13];
        Psram_Valid_To_Systolic_FIFO_14[12] <= Psram_Valid_To_Systolic_FIFO_14[13];
        Psram_Valid_To_Systolic_FIFO_15[12] <= Psram_Valid_To_Systolic_FIFO_15[13];
        Psram_Valid_To_Systolic_FIFO_16[12] <= Psram_Valid_To_Systolic_FIFO_16[13];
        Psram_Valid_To_Systolic_FIFO_17[12] <= Psram_Valid_To_Systolic_FIFO_17[13];
        Psram_Valid_To_Systolic_FIFO_18[12] <= Psram_Valid_To_Systolic_FIFO_18[13];
        Psram_Valid_To_Systolic_FIFO_19[12] <= Psram_Valid_To_Systolic_FIFO_19[13];
        Psram_Valid_To_Systolic_FIFO_20[12] <= Psram_Valid_To_Systolic_FIFO_20[13];
        Psram_Valid_To_Systolic_FIFO_21[12] <= Psram_Valid_To_Systolic_FIFO_21[13];
        Psram_Valid_To_Systolic_FIFO_22[12] <= Psram_Valid_To_Systolic_FIFO_22[13];
        Psram_Valid_To_Systolic_FIFO_23[12] <= Psram_Valid_To_Systolic_FIFO_23[13];
        Psram_Valid_To_Systolic_FIFO_24[12] <= Psram_Valid_To_Systolic_FIFO_24[13];
        Psram_Valid_To_Systolic_FIFO_25[12] <= Psram_Valid_To_Systolic_FIFO_25[13];
        Psram_Valid_To_Systolic_FIFO_26[12] <= Psram_Valid_To_Systolic_FIFO_26[13];
        Psram_Valid_To_Systolic_FIFO_27[12] <= Psram_Valid_To_Systolic_FIFO_27[13];
        Psram_Valid_To_Systolic_FIFO_28[12] <= Psram_Valid_To_Systolic_FIFO_28[13];
        Psram_Valid_To_Systolic_FIFO_29[12] <= Psram_Valid_To_Systolic_FIFO_29[13];
        Psram_Valid_To_Systolic_FIFO_30[12] <= Psram_Valid_To_Systolic_FIFO_30[13];
        Psram_Valid_To_Systolic_FIFO_31[12] <= Psram_Valid_To_Systolic_FIFO_31[13];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_14[13] <= i_Psram_Valid_1buf[14];
        Psram_Valid_To_Systolic_FIFO_15[13] <= Psram_Valid_To_Systolic_FIFO_15[14];
        Psram_Valid_To_Systolic_FIFO_16[13] <= Psram_Valid_To_Systolic_FIFO_16[14];
        Psram_Valid_To_Systolic_FIFO_17[13] <= Psram_Valid_To_Systolic_FIFO_17[14];
        Psram_Valid_To_Systolic_FIFO_18[13] <= Psram_Valid_To_Systolic_FIFO_18[14];
        Psram_Valid_To_Systolic_FIFO_19[13] <= Psram_Valid_To_Systolic_FIFO_19[14];
        Psram_Valid_To_Systolic_FIFO_20[13] <= Psram_Valid_To_Systolic_FIFO_20[14];
        Psram_Valid_To_Systolic_FIFO_21[13] <= Psram_Valid_To_Systolic_FIFO_21[14];
        Psram_Valid_To_Systolic_FIFO_22[13] <= Psram_Valid_To_Systolic_FIFO_22[14];
        Psram_Valid_To_Systolic_FIFO_23[13] <= Psram_Valid_To_Systolic_FIFO_23[14];
        Psram_Valid_To_Systolic_FIFO_24[13] <= Psram_Valid_To_Systolic_FIFO_24[14];
        Psram_Valid_To_Systolic_FIFO_25[13] <= Psram_Valid_To_Systolic_FIFO_25[14];
        Psram_Valid_To_Systolic_FIFO_26[13] <= Psram_Valid_To_Systolic_FIFO_26[14];
        Psram_Valid_To_Systolic_FIFO_27[13] <= Psram_Valid_To_Systolic_FIFO_27[14];
        Psram_Valid_To_Systolic_FIFO_28[13] <= Psram_Valid_To_Systolic_FIFO_28[14];
        Psram_Valid_To_Systolic_FIFO_29[13] <= Psram_Valid_To_Systolic_FIFO_29[14];
        Psram_Valid_To_Systolic_FIFO_30[13] <= Psram_Valid_To_Systolic_FIFO_30[14];
        Psram_Valid_To_Systolic_FIFO_31[13] <= Psram_Valid_To_Systolic_FIFO_31[14];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_15[14] <= i_Psram_Valid_1buf[15];
        Psram_Valid_To_Systolic_FIFO_16[14] <= Psram_Valid_To_Systolic_FIFO_16[15];
        Psram_Valid_To_Systolic_FIFO_17[14] <= Psram_Valid_To_Systolic_FIFO_17[15];
        Psram_Valid_To_Systolic_FIFO_18[14] <= Psram_Valid_To_Systolic_FIFO_18[15];
        Psram_Valid_To_Systolic_FIFO_19[14] <= Psram_Valid_To_Systolic_FIFO_19[15];
        Psram_Valid_To_Systolic_FIFO_20[14] <= Psram_Valid_To_Systolic_FIFO_20[15];
        Psram_Valid_To_Systolic_FIFO_21[14] <= Psram_Valid_To_Systolic_FIFO_21[15];
        Psram_Valid_To_Systolic_FIFO_22[14] <= Psram_Valid_To_Systolic_FIFO_22[15];
        Psram_Valid_To_Systolic_FIFO_23[14] <= Psram_Valid_To_Systolic_FIFO_23[15];
        Psram_Valid_To_Systolic_FIFO_24[14] <= Psram_Valid_To_Systolic_FIFO_24[15];
        Psram_Valid_To_Systolic_FIFO_25[14] <= Psram_Valid_To_Systolic_FIFO_25[15];
        Psram_Valid_To_Systolic_FIFO_26[14] <= Psram_Valid_To_Systolic_FIFO_26[15];
        Psram_Valid_To_Systolic_FIFO_27[14] <= Psram_Valid_To_Systolic_FIFO_27[15];
        Psram_Valid_To_Systolic_FIFO_28[14] <= Psram_Valid_To_Systolic_FIFO_28[15];
        Psram_Valid_To_Systolic_FIFO_29[14] <= Psram_Valid_To_Systolic_FIFO_29[15];
        Psram_Valid_To_Systolic_FIFO_30[14] <= Psram_Valid_To_Systolic_FIFO_30[15];
        Psram_Valid_To_Systolic_FIFO_31[14] <= Psram_Valid_To_Systolic_FIFO_31[15];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_16[15] <= i_Psram_Valid_1buf[16];
        Psram_Valid_To_Systolic_FIFO_17[15] <= Psram_Valid_To_Systolic_FIFO_17[16];
        Psram_Valid_To_Systolic_FIFO_18[15] <= Psram_Valid_To_Systolic_FIFO_18[16];
        Psram_Valid_To_Systolic_FIFO_19[15] <= Psram_Valid_To_Systolic_FIFO_19[16];
        Psram_Valid_To_Systolic_FIFO_20[15] <= Psram_Valid_To_Systolic_FIFO_20[16];
        Psram_Valid_To_Systolic_FIFO_21[15] <= Psram_Valid_To_Systolic_FIFO_21[16];
        Psram_Valid_To_Systolic_FIFO_22[15] <= Psram_Valid_To_Systolic_FIFO_22[16];
        Psram_Valid_To_Systolic_FIFO_23[15] <= Psram_Valid_To_Systolic_FIFO_23[16];
        Psram_Valid_To_Systolic_FIFO_24[15] <= Psram_Valid_To_Systolic_FIFO_24[16];
        Psram_Valid_To_Systolic_FIFO_25[15] <= Psram_Valid_To_Systolic_FIFO_25[16];
        Psram_Valid_To_Systolic_FIFO_26[15] <= Psram_Valid_To_Systolic_FIFO_26[16];
        Psram_Valid_To_Systolic_FIFO_27[15] <= Psram_Valid_To_Systolic_FIFO_27[16];
        Psram_Valid_To_Systolic_FIFO_28[15] <= Psram_Valid_To_Systolic_FIFO_28[16];
        Psram_Valid_To_Systolic_FIFO_29[15] <= Psram_Valid_To_Systolic_FIFO_29[16];
        Psram_Valid_To_Systolic_FIFO_30[15] <= Psram_Valid_To_Systolic_FIFO_30[16];
        Psram_Valid_To_Systolic_FIFO_31[15] <= Psram_Valid_To_Systolic_FIFO_31[16];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_17[16] <= i_Psram_Valid_1buf[17];
        Psram_Valid_To_Systolic_FIFO_18[16] <= Psram_Valid_To_Systolic_FIFO_18[17];
        Psram_Valid_To_Systolic_FIFO_19[16] <= Psram_Valid_To_Systolic_FIFO_19[17];
        Psram_Valid_To_Systolic_FIFO_20[16] <= Psram_Valid_To_Systolic_FIFO_20[17];
        Psram_Valid_To_Systolic_FIFO_21[16] <= Psram_Valid_To_Systolic_FIFO_21[17];
        Psram_Valid_To_Systolic_FIFO_22[16] <= Psram_Valid_To_Systolic_FIFO_22[17];
        Psram_Valid_To_Systolic_FIFO_23[16] <= Psram_Valid_To_Systolic_FIFO_23[17];
        Psram_Valid_To_Systolic_FIFO_24[16] <= Psram_Valid_To_Systolic_FIFO_24[17];
        Psram_Valid_To_Systolic_FIFO_25[16] <= Psram_Valid_To_Systolic_FIFO_25[17];
        Psram_Valid_To_Systolic_FIFO_26[16] <= Psram_Valid_To_Systolic_FIFO_26[17];
        Psram_Valid_To_Systolic_FIFO_27[16] <= Psram_Valid_To_Systolic_FIFO_27[17];
        Psram_Valid_To_Systolic_FIFO_28[16] <= Psram_Valid_To_Systolic_FIFO_28[17];
        Psram_Valid_To_Systolic_FIFO_29[16] <= Psram_Valid_To_Systolic_FIFO_29[17];
        Psram_Valid_To_Systolic_FIFO_30[16] <= Psram_Valid_To_Systolic_FIFO_30[17];
        Psram_Valid_To_Systolic_FIFO_31[16] <= Psram_Valid_To_Systolic_FIFO_31[17];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_18[17] <= i_Psram_Valid_1buf[18];
        Psram_Valid_To_Systolic_FIFO_19[17] <= Psram_Valid_To_Systolic_FIFO_19[18];
        Psram_Valid_To_Systolic_FIFO_20[17] <= Psram_Valid_To_Systolic_FIFO_20[18];
        Psram_Valid_To_Systolic_FIFO_21[17] <= Psram_Valid_To_Systolic_FIFO_21[18];
        Psram_Valid_To_Systolic_FIFO_22[17] <= Psram_Valid_To_Systolic_FIFO_22[18];
        Psram_Valid_To_Systolic_FIFO_23[17] <= Psram_Valid_To_Systolic_FIFO_23[18];
        Psram_Valid_To_Systolic_FIFO_24[17] <= Psram_Valid_To_Systolic_FIFO_24[18];
        Psram_Valid_To_Systolic_FIFO_25[17] <= Psram_Valid_To_Systolic_FIFO_25[18];
        Psram_Valid_To_Systolic_FIFO_26[17] <= Psram_Valid_To_Systolic_FIFO_26[18];
        Psram_Valid_To_Systolic_FIFO_27[17] <= Psram_Valid_To_Systolic_FIFO_27[18];
        Psram_Valid_To_Systolic_FIFO_28[17] <= Psram_Valid_To_Systolic_FIFO_28[18];
        Psram_Valid_To_Systolic_FIFO_29[17] <= Psram_Valid_To_Systolic_FIFO_29[18];
        Psram_Valid_To_Systolic_FIFO_30[17] <= Psram_Valid_To_Systolic_FIFO_30[18];
        Psram_Valid_To_Systolic_FIFO_31[17] <= Psram_Valid_To_Systolic_FIFO_31[18];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_19[18] <= i_Psram_Valid_1buf[19];
        Psram_Valid_To_Systolic_FIFO_20[18] <= Psram_Valid_To_Systolic_FIFO_20[19];
        Psram_Valid_To_Systolic_FIFO_21[18] <= Psram_Valid_To_Systolic_FIFO_21[19];
        Psram_Valid_To_Systolic_FIFO_22[18] <= Psram_Valid_To_Systolic_FIFO_22[19];
        Psram_Valid_To_Systolic_FIFO_23[18] <= Psram_Valid_To_Systolic_FIFO_23[19];
        Psram_Valid_To_Systolic_FIFO_24[18] <= Psram_Valid_To_Systolic_FIFO_24[19];
        Psram_Valid_To_Systolic_FIFO_25[18] <= Psram_Valid_To_Systolic_FIFO_25[19];
        Psram_Valid_To_Systolic_FIFO_26[18] <= Psram_Valid_To_Systolic_FIFO_26[19];
        Psram_Valid_To_Systolic_FIFO_27[18] <= Psram_Valid_To_Systolic_FIFO_27[19];
        Psram_Valid_To_Systolic_FIFO_28[18] <= Psram_Valid_To_Systolic_FIFO_28[19];
        Psram_Valid_To_Systolic_FIFO_29[18] <= Psram_Valid_To_Systolic_FIFO_29[19];
        Psram_Valid_To_Systolic_FIFO_30[18] <= Psram_Valid_To_Systolic_FIFO_30[19];
        Psram_Valid_To_Systolic_FIFO_31[18] <= Psram_Valid_To_Systolic_FIFO_31[19];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_20[19] <= i_Psram_Valid_1buf[20];
        Psram_Valid_To_Systolic_FIFO_21[19] <= Psram_Valid_To_Systolic_FIFO_21[20];
        Psram_Valid_To_Systolic_FIFO_22[19] <= Psram_Valid_To_Systolic_FIFO_22[20];
        Psram_Valid_To_Systolic_FIFO_23[19] <= Psram_Valid_To_Systolic_FIFO_23[20];
        Psram_Valid_To_Systolic_FIFO_24[19] <= Psram_Valid_To_Systolic_FIFO_24[20];
        Psram_Valid_To_Systolic_FIFO_25[19] <= Psram_Valid_To_Systolic_FIFO_25[20];
        Psram_Valid_To_Systolic_FIFO_26[19] <= Psram_Valid_To_Systolic_FIFO_26[20];
        Psram_Valid_To_Systolic_FIFO_27[19] <= Psram_Valid_To_Systolic_FIFO_27[20];
        Psram_Valid_To_Systolic_FIFO_28[19] <= Psram_Valid_To_Systolic_FIFO_28[20];
        Psram_Valid_To_Systolic_FIFO_29[19] <= Psram_Valid_To_Systolic_FIFO_29[20];
        Psram_Valid_To_Systolic_FIFO_30[19] <= Psram_Valid_To_Systolic_FIFO_30[20];
        Psram_Valid_To_Systolic_FIFO_31[19] <= Psram_Valid_To_Systolic_FIFO_31[20];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_21[20] <= i_Psram_Valid_1buf[21];
        Psram_Valid_To_Systolic_FIFO_22[20] <= Psram_Valid_To_Systolic_FIFO_22[21];
        Psram_Valid_To_Systolic_FIFO_23[20] <= Psram_Valid_To_Systolic_FIFO_23[21];
        Psram_Valid_To_Systolic_FIFO_24[20] <= Psram_Valid_To_Systolic_FIFO_24[21];
        Psram_Valid_To_Systolic_FIFO_25[20] <= Psram_Valid_To_Systolic_FIFO_25[21];
        Psram_Valid_To_Systolic_FIFO_26[20] <= Psram_Valid_To_Systolic_FIFO_26[21];
        Psram_Valid_To_Systolic_FIFO_27[20] <= Psram_Valid_To_Systolic_FIFO_27[21];
        Psram_Valid_To_Systolic_FIFO_28[20] <= Psram_Valid_To_Systolic_FIFO_28[21];
        Psram_Valid_To_Systolic_FIFO_29[20] <= Psram_Valid_To_Systolic_FIFO_29[21];
        Psram_Valid_To_Systolic_FIFO_30[20] <= Psram_Valid_To_Systolic_FIFO_30[21];
        Psram_Valid_To_Systolic_FIFO_31[20] <= Psram_Valid_To_Systolic_FIFO_31[21];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_22[21] <= i_Psram_Valid_1buf[22];
        Psram_Valid_To_Systolic_FIFO_23[21] <= Psram_Valid_To_Systolic_FIFO_23[22];
        Psram_Valid_To_Systolic_FIFO_24[21] <= Psram_Valid_To_Systolic_FIFO_24[22];
        Psram_Valid_To_Systolic_FIFO_25[21] <= Psram_Valid_To_Systolic_FIFO_25[22];
        Psram_Valid_To_Systolic_FIFO_26[21] <= Psram_Valid_To_Systolic_FIFO_26[22];
        Psram_Valid_To_Systolic_FIFO_27[21] <= Psram_Valid_To_Systolic_FIFO_27[22];
        Psram_Valid_To_Systolic_FIFO_28[21] <= Psram_Valid_To_Systolic_FIFO_28[22];
        Psram_Valid_To_Systolic_FIFO_29[21] <= Psram_Valid_To_Systolic_FIFO_29[22];
        Psram_Valid_To_Systolic_FIFO_30[21] <= Psram_Valid_To_Systolic_FIFO_30[22];
        Psram_Valid_To_Systolic_FIFO_31[21] <= Psram_Valid_To_Systolic_FIFO_31[22];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_23[22] <= i_Psram_Valid_1buf[23];
        Psram_Valid_To_Systolic_FIFO_24[22] <= Psram_Valid_To_Systolic_FIFO_24[23];
        Psram_Valid_To_Systolic_FIFO_25[22] <= Psram_Valid_To_Systolic_FIFO_25[23];
        Psram_Valid_To_Systolic_FIFO_26[22] <= Psram_Valid_To_Systolic_FIFO_26[23];
        Psram_Valid_To_Systolic_FIFO_27[22] <= Psram_Valid_To_Systolic_FIFO_27[23];
        Psram_Valid_To_Systolic_FIFO_28[22] <= Psram_Valid_To_Systolic_FIFO_28[23];
        Psram_Valid_To_Systolic_FIFO_29[22] <= Psram_Valid_To_Systolic_FIFO_29[23];
        Psram_Valid_To_Systolic_FIFO_30[22] <= Psram_Valid_To_Systolic_FIFO_30[23];
        Psram_Valid_To_Systolic_FIFO_31[22] <= Psram_Valid_To_Systolic_FIFO_31[23];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_24[23] <= i_Psram_Valid_1buf[24];
        Psram_Valid_To_Systolic_FIFO_25[23] <= Psram_Valid_To_Systolic_FIFO_25[24];
        Psram_Valid_To_Systolic_FIFO_26[23] <= Psram_Valid_To_Systolic_FIFO_26[24];
        Psram_Valid_To_Systolic_FIFO_27[23] <= Psram_Valid_To_Systolic_FIFO_27[24];
        Psram_Valid_To_Systolic_FIFO_28[23] <= Psram_Valid_To_Systolic_FIFO_28[24];
        Psram_Valid_To_Systolic_FIFO_29[23] <= Psram_Valid_To_Systolic_FIFO_29[24];
        Psram_Valid_To_Systolic_FIFO_30[23] <= Psram_Valid_To_Systolic_FIFO_30[24];
        Psram_Valid_To_Systolic_FIFO_31[23] <= Psram_Valid_To_Systolic_FIFO_31[24];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_25[24] <= i_Psram_Valid_1buf[25];
        Psram_Valid_To_Systolic_FIFO_26[24] <= Psram_Valid_To_Systolic_FIFO_26[25];
        Psram_Valid_To_Systolic_FIFO_27[24] <= Psram_Valid_To_Systolic_FIFO_27[25];
        Psram_Valid_To_Systolic_FIFO_28[24] <= Psram_Valid_To_Systolic_FIFO_28[25];
        Psram_Valid_To_Systolic_FIFO_29[24] <= Psram_Valid_To_Systolic_FIFO_29[25];
        Psram_Valid_To_Systolic_FIFO_30[24] <= Psram_Valid_To_Systolic_FIFO_30[25];
        Psram_Valid_To_Systolic_FIFO_31[24] <= Psram_Valid_To_Systolic_FIFO_31[25];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_26[25] <= i_Psram_Valid_1buf[26];
        Psram_Valid_To_Systolic_FIFO_27[25] <= Psram_Valid_To_Systolic_FIFO_27[26];
        Psram_Valid_To_Systolic_FIFO_28[25] <= Psram_Valid_To_Systolic_FIFO_28[26];
        Psram_Valid_To_Systolic_FIFO_29[25] <= Psram_Valid_To_Systolic_FIFO_29[26];
        Psram_Valid_To_Systolic_FIFO_30[25] <= Psram_Valid_To_Systolic_FIFO_30[26];
        Psram_Valid_To_Systolic_FIFO_31[25] <= Psram_Valid_To_Systolic_FIFO_31[26];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_27[26] <= i_Psram_Valid_1buf[27];
        Psram_Valid_To_Systolic_FIFO_28[26] <= Psram_Valid_To_Systolic_FIFO_28[27];
        Psram_Valid_To_Systolic_FIFO_29[26] <= Psram_Valid_To_Systolic_FIFO_29[27];
        Psram_Valid_To_Systolic_FIFO_30[26] <= Psram_Valid_To_Systolic_FIFO_30[27];
        Psram_Valid_To_Systolic_FIFO_31[26] <= Psram_Valid_To_Systolic_FIFO_31[27];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_28[27] <= i_Psram_Valid_1buf[28];
        Psram_Valid_To_Systolic_FIFO_29[27] <= Psram_Valid_To_Systolic_FIFO_29[28];
        Psram_Valid_To_Systolic_FIFO_30[27] <= Psram_Valid_To_Systolic_FIFO_30[28];
        Psram_Valid_To_Systolic_FIFO_31[27] <= Psram_Valid_To_Systolic_FIFO_31[28];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_29[28] <= i_Psram_Valid_1buf[29];
        Psram_Valid_To_Systolic_FIFO_30[28] <= Psram_Valid_To_Systolic_FIFO_30[29];
        Psram_Valid_To_Systolic_FIFO_31[28] <= Psram_Valid_To_Systolic_FIFO_31[29];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_30[29] <= i_Psram_Valid_1buf[30];
        Psram_Valid_To_Systolic_FIFO_31[29] <= Psram_Valid_To_Systolic_FIFO_31[30];
    end

    always @(posedge CLK) begin
        Psram_Valid_To_Systolic_FIFO_31[30] <= i_Psram_Valid_1buf[31];
    end

endmodule